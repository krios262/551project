module VADD(arguments)

endmodule
