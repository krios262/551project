module SMUL16(output reg [255:0] product,output reg Ovf, input [15:0] scalar,input [255:0] vecin);

SMUL(product[255:240],Ovf,scalar[15:0], vecin[255:240]);
SMUL(product[239:224],Ovf,scalar[15:0], vecin[239:224]);
SMUL(product[223:208],Ovf,scalar[15:0], vecin[223:208]);
SMUL(product[207:192],Ovf,scalar[15:0], vecin[207:192]);
SMUL(product[191:176],Ovf,scalar[15:0], vecin[191:176]);
SMUL(product[175:160],Ovf,scalar[15:0], vecin[175:160]);
SMUL(product[159:144],Ovf,scalar[15:0], vecin[159:144]);
SMUL(product[143:128],Ovf,scalar[15:0], vecin[143:128]);
SMUL(product[127:112],Ovf,scalar[15:0], vecin[127:112]);
SMUL(product[111:96],Ovf,scalar[15:0], vecin[111:96]);
SMUL(product[95:80],Ovf,scalar[15:0], vecin[95:80]);
SMUL(product[79:64],Ovf,scalar[15:0], vecin[79:64]);
SMUL(product[63:48],Ovf,scalar[15:0], vecin[63:48]);
SMUL(product[47:32],Ovf,scalar[15:0], vecin[47:32]);
SMUL(product[31:16],Ovf,scalar[15:0], vecin[31:16]);
SMUL(product[15:0],Ovf,scalar[15:0], vecin[15:0]);

endmodule

module t_SMULv();
  
  wire [255:0] pro;
  
  reg [255:0] vec1;
  reg [15:0] s1;
  
  SMUL16 S1(pro,s1,vec1);
  
  initial begin
    s1 = 16'hA;
    vec1 = 256'h00010203;
    #10 vec1 = 256'h00020304;
    #20 vec1 = 256'h0406080a;
end
endmodule

module SMUL(output reg [15:0] prod,output reg Overflow,input [15:0] A, input [15:0] B, output reg [22:0] operprod,output reg [6:0] temp_exp);
  
  reg [11:0] operA,operB;
  wire [11:0] operA1,operB1,operA2,operB2;
  //reg [23:0] operprod;
  reg [9:0] operprod1;
  reg [11:0] operprod2;
  reg [5:0] i = 6'b000000;
  reg [5:0] j = 4'b0000;
  reg [1:0] oper;
  reg flag;
  reg flagz;
  //reg [6:0] temp_exp;
  
  //append sticky and guard bit along with normalised one
  assign operA1 = {1'b0,1'b1,A[9:0]};
  assign operB1 = {1'b0,1'b1,B[9:0]}; 
  assign operA2 = {2'b0,A[9:0]};
  assign operB2 = {2'b0,B[9:0]};
  
  //perform floating point multiplication
  always @(*)
  //check if any number is infinity if so make the product equal to infinity
  begin
  if((A[14:10] == 5'h1F) || (B[14:10] == 5'h1F))
  begin
     if (A[14:10] == 5'h1F) 
       begin
         prod = {A[15],A[14:10],10'h0};
         Overflow = 1'b1;
       end
     else 
       begin
         prod = {B[15],B[14:10],10'h0};
         Overflow = 1'b1;
       end
  end
  //based on whether the number is normalised or denormalised build the inputs for the multiplication
  else
  begin
  if((A[14:10] == 5'h0) && (B[14:10] == 5'h0))
  begin 
    operA = operA2;
    operB = operB2;
  end
  else if (A[14:10] == 5'h0)
  begin
    operA = operA2;
    operB = operB1;
  end
  else if(B[14:10] == 5'h0)
  begin
    operA = operA1;
    operB = operB2;
  end
  else
  begin
    operA = operA1;
    operB = operB1;
  end
  
  //calculate temp exponent
  temp_exp = A[14:10]+B[14:10]- 4'hf;
  
  //calculate the product of two 11 bit numbers
  operprod = operA*operB;
  
  
  // if temp_exp is greater than 31 it is a denormalised number
  if (temp_exp > 5'h1e)
    begin
       prod[15] = A[15] ^ B[15];
       prod[14:10] = 5'd31;
       prod[9:0] = 10'h0;
    end
    
  // if the last bit is set do the following
  else
    begin
    if(operprod[21] == 1'b1)
    begin
    if (temp_exp > 5'h1d)
      begin
        prod[15] = A[15] ^ B[15];
        prod[14:10] = 5'd31;
        prod[9:0] = 10'h0;
      end
    else
      begin
        prod[15] = A[15] ^ B[15];
        //rounding off logic
          if(operprod[10] == 1'b1 && operprod[11] == 1'b1)
            begin
              operprod2 = operprod[21:11]+1;
            end
          else
            begin
              operprod2 = operprod[21:11];
            end
          // exponent reassign and normalise after rounding
          if(operprod2[11] == 1'b1 && temp_exp < 5'h1d)
            begin
              prod[14:10] = temp_exp+2;
              operprod1[9:0] = operprod2[10:1];
              Overflow = 1'b0;
            end
           else if((operprod2[11] == 1'b1 && temp_exp == 5'h1d)||(operprod2[10] == 1'b1 && temp_exp == 5'h1e))
            begin
              prod[14:10] = 5'd31;
              operprod1[9:0] = 10'h1;
              Overflow = 1'b0;
            end         
           else        
            begin
              prod[14:10] = temp_exp+1;
              operprod1[9:0] = operprod2[9:0];
              Overflow = 1'b0;
            end 
          end
        end
        
     // if 21st bit of product is 1
     else if(operprod[20] == 1'b1)
      begin
        prod[15] = A[15] ^ B[15];
        //rounding off logic
          if(operprod[10] == 1'b1 && operprod[9] == 1'b1)
            begin
              operprod2 = operprod[19:10]+1;
            end
          else
            begin
              operprod2 = operprod[19:10];
            end
          // exponent reassign and normalise after rounding
          if(operprod2[11] == 1'b1 && temp_exp < 5'h1e)
            begin
              prod[14:10] = temp_exp+1;
              Overflow = 1'b0;
              operprod1[9:0] = operprod2[10:1];
            end
           else if(operprod2[11] == 1'b1 && temp_exp == 5'h1e)
            begin
              prod[14:10] = 5'd31;
              Overflow = 1'b1;
              operprod1[9:0] = 10'h0;
            end
          else
            begin
              prod[14:10] = temp_exp;
              operprod1[9:0] = operprod2[9:0];
              Overflow = 1'b0;
            end
          end
          
    // if a denormalised number is a part of input for multiplication
    else
      begin
        flag =1'b0;
        flagz = 1'b0;
        Overflow = 1'b0;
        for(j=0;j<22;j=j+1)
          begin
            if(((operprod[20])== 1'b0))
              begin
                if((flag == 1'b0) && (flagz == 1'b0))
                  begin
                    operprod = operprod << 1'b1;
                    temp_exp = temp_exp - 1'b1; 
                    if(temp_exp == 1'b0)
                      begin
                        flagz = 1'b1;
                      end
                    else
                      begin
                        flagz = 1'b0;
                      end
                  end
                end
            else
              begin
                operprod = operprod;
                temp_exp = temp_exp;
                flag = 1'b1;
              end
         end
         
         if((operprod[20] ==  1'b1) && (temp_exp ==7'b0))
           begin
             temp_exp= temp_exp+1'b1;
           end
         else
           begin
             temp_exp = temp_exp;
           end
         
            // calculating the sign
           prod[15] = A[15] ^ B[15];
           //rounding off logic
          if(operprod[10] == 1'b1 && operprod[9] == 1'b1)
            begin
              operprod2 = operprod[19:10]+1;
            end
          else
            begin
              operprod2 = operprod[19:10];
            end
          // exponent reassign and normalise after rounding
          if(operprod2[11] == 1'b1 && temp_exp < 5'h1e)
            begin
              prod[14:10] = temp_exp+1;
              Overflow = 1'b0;
              operprod1[9:0] = operprod2[10:1];
            end
          else
            begin
              prod[14:10] = temp_exp;
              operprod1[9:0] = operprod2[9:0];
              Overflow = 1'b0;
            end
       end
      prod[9:0] = operprod1;
        
      end  
      end
    end
    endmodule
            
            
module t_SMUL();
  
  wire [15:0] prd;
  wire ov;
  wire [6:0] ex;
  reg [15:0] vect;
  reg [15:0] sa;
  wire [22:0] mant;
  
  SMUL S1(prd,ov,sa,vect,mant,ex);
  
  initial begin
    sa = 16'h4080;
    vect = 16'h0011;
    
    #20 sa = 16'h4080;
    vect = 16'h0201;
    
end
endmodule            
      
`timescale 100ps/1ps
module t_SMUL_synth();
  
  wire [15:0] prd;
  wire ov;
  wire [6:0] ex;
  reg [15:0] vect;
  reg [15:0] sa;
  wire [22:0] mant;
  
  SMUL_synth S1(prd,ov,sa,vect,mant,ex);
  
  initial begin
    sa = 16'h4080;
    vect = 16'h0011;
    
    #20 sa = 16'h4080;
    vect = 16'h0201;
    
end
endmodule 
 

module SMUL_synth ( prod, Overflow, A, B, operprod, temp_exp );
  output [15:0] prod;
  input [15:0] A;
  input [15:0] B;
  output [22:0] operprod;
  output [6:0] temp_exp;
  output Overflow;
  wire   N78, N92, N93, N107, N108, N109, N110, N111, N112, N113, N114, N115,
         N116, N117, N118, N119, N120, N121, N122, N123, N124, N125, N126,
         N127, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N1782, N1783, N1784, N1785, N1786, N1787, N1788, N1789, N1790, N1791,
         N1846, N1847, N1848, N1849, N1850, N1851, N1852, N1853, N1854, N1855,
         N1911, N1912, N1913, N1914, N1915, N1916, N1917, N1919, N1920, N1921,
         N1922, N1923, N1924, N1925, N1926, N1927, N1928, N1929, N1930, N1931,
         N1932, N1933, N1934, N1935, N1936, N1937, N1938, N1939, N1940, N1942,
         \C148/DATA4_0 , \C148/DATA4_1 , \C148/DATA4_2 , \C148/DATA4_3 ,
         \C148/DATA4_4 , \C148/DATA4_5 , \C148/DATA4_6 , \C148/DATA4_7 ,
         \C148/DATA4_8 , \DP_OP_379J1_125_371/I4 , \DP_OP_379J1_125_371/I5 ,
         \DP_OP_379J1_125_371/n342 , \DP_OP_379J1_125_371/n341 ,
         \DP_OP_379J1_125_371/n340 , \DP_OP_379J1_125_371/n339 ,
         \DP_OP_379J1_125_371/n338 , \DP_OP_379J1_125_371/n337 ,
         \DP_OP_379J1_125_371/n336 , \DP_OP_379J1_125_371/n335 ,
         \DP_OP_379J1_125_371/n329 , \DP_OP_379J1_125_371/n328 ,
         \DP_OP_379J1_125_371/n327 , \DP_OP_379J1_125_371/n326 ,
         \DP_OP_379J1_125_371/n325 , \DP_OP_379J1_125_371/n324 ,
         \DP_OP_379J1_125_371/n323 , \DP_OP_379J1_125_371/n322 ,
         \DP_OP_379J1_125_371/n321 , \DP_OP_379J1_125_371/n320 ,
         \DP_OP_379J1_125_371/n319 , \DP_OP_379J1_125_371/n279 ,
         \DP_OP_379J1_125_371/n278 , \DP_OP_379J1_125_371/n277 ,
         \DP_OP_379J1_125_371/n276 , \DP_OP_379J1_125_371/n275 ,
         \DP_OP_379J1_125_371/n274 , \DP_OP_379J1_125_371/n273 ,
         \DP_OP_379J1_125_371/n272 , \DP_OP_379J1_125_371/n271 ,
         \DP_OP_379J1_125_371/n270 , \DP_OP_379J1_125_371/n269 ,
         \DP_OP_379J1_125_371/n268 , \DP_OP_379J1_125_371/n267 ,
         \DP_OP_379J1_125_371/n266 , \DP_OP_379J1_125_371/n265 ,
         \DP_OP_379J1_125_371/n264 , \DP_OP_379J1_125_371/n263 ,
         \DP_OP_379J1_125_371/n262 , \DP_OP_379J1_125_371/n261 ,
         \DP_OP_379J1_125_371/n260 , \DP_OP_379J1_125_371/n259 ,
         \DP_OP_379J1_125_371/n258 , \DP_OP_379J1_125_371/n257 ,
         \DP_OP_379J1_125_371/n256 , \DP_OP_379J1_125_371/n255 ,
         \DP_OP_379J1_125_371/n254 , \DP_OP_379J1_125_371/n253 ,
         \DP_OP_379J1_125_371/n252 , \DP_OP_379J1_125_371/n251 ,
         \DP_OP_379J1_125_371/n250 , \DP_OP_379J1_125_371/n249 ,
         \DP_OP_379J1_125_371/n248 , \DP_OP_379J1_125_371/n247 ,
         \DP_OP_379J1_125_371/n246 , \DP_OP_379J1_125_371/n245 ,
         \DP_OP_379J1_125_371/n244 , \DP_OP_379J1_125_371/n243 ,
         \DP_OP_379J1_125_371/n242 , \DP_OP_379J1_125_371/n241 ,
         \DP_OP_379J1_125_371/n240 , \DP_OP_379J1_125_371/n239 ,
         \DP_OP_379J1_125_371/n238 , \DP_OP_379J1_125_371/n237 ,
         \DP_OP_379J1_125_371/n236 , \DP_OP_379J1_125_371/n235 ,
         \DP_OP_379J1_125_371/n234 , \DP_OP_379J1_125_371/n233 ,
         \DP_OP_379J1_125_371/n232 , \DP_OP_379J1_125_371/n231 ,
         \DP_OP_379J1_125_371/n230 , \DP_OP_379J1_125_371/n229 ,
         \DP_OP_379J1_125_371/n228 , \DP_OP_379J1_125_371/n227 ,
         \DP_OP_379J1_125_371/n226 , \DP_OP_379J1_125_371/n225 ,
         \DP_OP_379J1_125_371/n224 , \DP_OP_379J1_125_371/n223 ,
         \DP_OP_379J1_125_371/n222 , \DP_OP_379J1_125_371/n221 ,
         \DP_OP_379J1_125_371/n220 , \DP_OP_379J1_125_371/n208 ,
         \DP_OP_379J1_125_371/n207 , \DP_OP_379J1_125_371/n206 ,
         \DP_OP_379J1_125_371/n205 , \DP_OP_379J1_125_371/n204 ,
         \DP_OP_379J1_125_371/n203 , \DP_OP_379J1_125_371/n202 ,
         \DP_OP_379J1_125_371/n201 , \DP_OP_379J1_125_371/n200 ,
         \DP_OP_379J1_125_371/n199 , \DP_OP_379J1_125_371/n198 ,
         \DP_OP_379J1_125_371/n197 , \DP_OP_379J1_125_371/n196 ,
         \DP_OP_379J1_125_371/n195 , \DP_OP_379J1_125_371/n194 ,
         \DP_OP_379J1_125_371/n193 , \DP_OP_379J1_125_371/n192 ,
         \DP_OP_379J1_125_371/n191 , \DP_OP_379J1_125_371/n190 ,
         \DP_OP_379J1_125_371/n189 , \DP_OP_379J1_125_371/n188 ,
         \DP_OP_379J1_125_371/n187 , \DP_OP_379J1_125_371/n186 ,
         \DP_OP_379J1_125_371/n185 , \DP_OP_379J1_125_371/n184 ,
         \DP_OP_379J1_125_371/n183 , \DP_OP_379J1_125_371/n182 ,
         \DP_OP_379J1_125_371/n181 , \DP_OP_379J1_125_371/n180 ,
         \DP_OP_379J1_125_371/n179 , \DP_OP_379J1_125_371/n178 ,
         \DP_OP_379J1_125_371/n177 , \DP_OP_379J1_125_371/n176 ,
         \DP_OP_379J1_125_371/n175 , \DP_OP_379J1_125_371/n174 ,
         \DP_OP_379J1_125_371/n173 , \DP_OP_379J1_125_371/n172 ,
         \DP_OP_379J1_125_371/n171 , \DP_OP_379J1_125_371/n170 ,
         \DP_OP_379J1_125_371/n169 , \DP_OP_379J1_125_371/n168 ,
         \DP_OP_379J1_125_371/n167 , \DP_OP_379J1_125_371/n166 ,
         \DP_OP_379J1_125_371/n165 , \DP_OP_379J1_125_371/n164 ,
         \DP_OP_379J1_125_371/n163 , \DP_OP_379J1_125_371/n162 ,
         \DP_OP_379J1_125_371/n161 , \DP_OP_379J1_125_371/n160 ,
         \DP_OP_379J1_125_371/n159 , \DP_OP_379J1_125_371/n158 ,
         \DP_OP_379J1_125_371/n157 , \DP_OP_379J1_125_371/n156 ,
         \DP_OP_379J1_125_371/n155 , \DP_OP_379J1_125_371/n154 ,
         \DP_OP_379J1_125_371/n153 , \DP_OP_379J1_125_371/n152 ,
         \DP_OP_379J1_125_371/n151 , \DP_OP_379J1_125_371/n150 ,
         \DP_OP_379J1_125_371/n149 , \DP_OP_379J1_125_371/n148 ,
         \DP_OP_379J1_125_371/n147 , \DP_OP_379J1_125_371/n146 ,
         \DP_OP_379J1_125_371/n145 , \DP_OP_379J1_125_371/n144 ,
         \DP_OP_379J1_125_371/n143 , \DP_OP_379J1_125_371/n142 ,
         \DP_OP_379J1_125_371/n141 , \DP_OP_379J1_125_371/n140 ,
         \DP_OP_379J1_125_371/n139 , \DP_OP_379J1_125_371/n138 ,
         \DP_OP_379J1_125_371/n136 , \DP_OP_379J1_125_371/n135 ,
         \DP_OP_379J1_125_371/n134 , \DP_OP_379J1_125_371/n133 ,
         \DP_OP_379J1_125_371/n132 , \DP_OP_379J1_125_371/n131 ,
         \DP_OP_379J1_125_371/n130 , \DP_OP_379J1_125_371/n129 ,
         \DP_OP_379J1_125_371/n128 , \DP_OP_379J1_125_371/n127 ,
         \DP_OP_379J1_125_371/n126 , \DP_OP_379J1_125_371/n125 ,
         \DP_OP_379J1_125_371/n124 , \DP_OP_379J1_125_371/n123 ,
         \DP_OP_379J1_125_371/n122 , \DP_OP_379J1_125_371/n121 ,
         \DP_OP_379J1_125_371/n120 , \DP_OP_379J1_125_371/n119 ,
         \DP_OP_379J1_125_371/n118 , \DP_OP_379J1_125_371/n117 ,
         \DP_OP_379J1_125_371/n116 , \DP_OP_379J1_125_371/n115 ,
         \DP_OP_379J1_125_371/n114 , \DP_OP_379J1_125_371/n113 ,
         \DP_OP_379J1_125_371/n112 , \DP_OP_379J1_125_371/n111 ,
         \DP_OP_379J1_125_371/n110 , \DP_OP_379J1_125_371/n109 ,
         \DP_OP_379J1_125_371/n108 , \DP_OP_379J1_125_371/n107 ,
         \DP_OP_379J1_125_371/n106 , \DP_OP_379J1_125_371/n105 ,
         \DP_OP_379J1_125_371/n104 , \DP_OP_379J1_125_371/n103 ,
         \DP_OP_379J1_125_371/n102 , \DP_OP_379J1_125_371/n101 ,
         \DP_OP_379J1_125_371/n100 , \DP_OP_379J1_125_371/n99 ,
         \DP_OP_379J1_125_371/n98 , \DP_OP_379J1_125_371/n97 ,
         \DP_OP_379J1_125_371/n96 , \DP_OP_379J1_125_371/n95 ,
         \DP_OP_379J1_125_371/n94 , \DP_OP_379J1_125_371/n93 ,
         \DP_OP_379J1_125_371/n92 , \DP_OP_379J1_125_371/n90 ,
         \DP_OP_379J1_125_371/n89 , \DP_OP_379J1_125_371/n88 ,
         \DP_OP_379J1_125_371/n87 , \DP_OP_379J1_125_371/n86 ,
         \DP_OP_379J1_125_371/n85 , \DP_OP_379J1_125_371/n83 ,
         \DP_OP_379J1_125_371/n82 , \DP_OP_379J1_125_371/n81 ,
         \DP_OP_379J1_125_371/n80 , \DP_OP_379J1_125_371/n79 ,
         \DP_OP_379J1_125_371/n78 , \DP_OP_379J1_125_371/n77 ,
         \DP_OP_379J1_125_371/n76 , \DP_OP_379J1_125_371/n75 ,
         \DP_OP_379J1_125_371/n74 , \DP_OP_379J1_125_371/n73 ,
         \DP_OP_379J1_125_371/n72 , \DP_OP_379J1_125_371/n71 ,
         \DP_OP_379J1_125_371/n69 , \DP_OP_379J1_125_371/n68 ,
         \DP_OP_379J1_125_371/n67 , \DP_OP_379J1_125_371/n66 ,
         \DP_OP_379J1_125_371/n65 , \DP_OP_379J1_125_371/n64 ,
         \DP_OP_379J1_125_371/n63 , \DP_OP_379J1_125_371/n62 ,
         \DP_OP_379J1_125_371/n61 , \DP_OP_379J1_125_371/n60 ,
         \DP_OP_379J1_125_371/n59 , \DP_OP_379J1_125_371/n57 ,
         \DP_OP_379J1_125_371/n56 , \DP_OP_379J1_125_371/n55 ,
         \DP_OP_379J1_125_371/n54 , \DP_OP_379J1_125_371/n53 ,
         \DP_OP_379J1_125_371/n52 , \DP_OP_379J1_125_371/n51 ,
         \DP_OP_379J1_125_371/n49 , \DP_OP_379J1_125_371/n48 ,
         \DP_OP_379J1_125_371/n47 , \DP_OP_379J1_125_371/n46 ,
         \DP_OP_379J1_125_371/n45 , \DP_OP_379J1_125_371/n43 ,
         \DP_OP_379J1_125_371/n42 , \DP_OP_379J1_125_371/n41 ,
         \DP_OP_379J1_125_371/n40 , \DP_OP_379J1_125_371/n39 ,
         \DP_OP_379J1_125_371/n38 , \DP_OP_379J1_125_371/n37 ,
         \DP_OP_379J1_125_371/n36 , \DP_OP_379J1_125_371/n35 ,
         \DP_OP_379J1_125_371/n34 , \DP_OP_379J1_125_371/n33 ,
         \DP_OP_379J1_125_371/n32 , \DP_OP_379J1_125_371/n31 ,
         \DP_OP_379J1_125_371/n30 , \DP_OP_379J1_125_371/n29 ,
         \DP_OP_379J1_125_371/n28 , \DP_OP_379J1_125_371/n27 ,
         \DP_OP_379J1_125_371/n26 , \DP_OP_379J1_125_371/n25 ,
         \DP_OP_379J1_125_371/n24 , \DP_OP_379J1_125_371/n19 ,
         \DP_OP_379J1_125_371/n18 , \DP_OP_379J1_125_371/n17 ,
         \DP_OP_379J1_125_371/n16 , \DP_OP_379J1_125_371/n15 ,
         \DP_OP_379J1_125_371/n14 , \DP_OP_379J1_125_371/n13 ,
         \DP_OP_379J1_125_371/n12 , \DP_OP_379J1_125_371/n11 ,
         \DP_OP_379J1_125_371/n10 , \DP_OP_379J1_125_371/n9 ,
         \DP_OP_379J1_125_371/n8 , \DP_OP_379J1_125_371/n7 ,
         \DP_OP_379J1_125_371/n6 , \DP_OP_379J1_125_371/n5 ,
         \DP_OP_379J1_125_371/n4 , \DP_OP_379J1_125_371/n3 ,
         \DP_OP_379J1_125_371/n2 , \DP_OP_379J1_125_371/n1 , n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350;
  wire   [9:0] operprod1;

  LNQD1BWP \operprod_reg[21]  ( .D(N1940), .EN(N78), .Q(operprod[21]) );
  LNQD1BWP \operprod_reg[20]  ( .D(N1939), .EN(N78), .Q(operprod[20]) );
  LNQD1BWP \operprod_reg[19]  ( .D(N1938), .EN(N78), .Q(operprod[19]) );
  LNQD1BWP \operprod_reg[18]  ( .D(N1937), .EN(N78), .Q(operprod[18]) );
  LNQD1BWP \operprod_reg[17]  ( .D(N1936), .EN(N78), .Q(operprod[17]) );
  LNQD1BWP \operprod_reg[16]  ( .D(N1935), .EN(N78), .Q(operprod[16]) );
  LNQD1BWP \operprod_reg[15]  ( .D(N1934), .EN(N78), .Q(operprod[15]) );
  LNQD1BWP \operprod_reg[14]  ( .D(N1933), .EN(N78), .Q(operprod[14]) );
  LNQD1BWP \operprod_reg[13]  ( .D(N1932), .EN(N78), .Q(operprod[13]) );
  LNQD1BWP \operprod_reg[12]  ( .D(N1931), .EN(N78), .Q(operprod[12]) );
  LNQD1BWP \operprod_reg[11]  ( .D(N1930), .EN(N78), .Q(operprod[11]) );
  LNQD1BWP \operprod_reg[10]  ( .D(N1929), .EN(N78), .Q(operprod[10]) );
  LNQD1BWP \operprod_reg[9]  ( .D(N1928), .EN(N78), .Q(operprod[9]) );
  LNQD1BWP \operprod_reg[8]  ( .D(N1927), .EN(N78), .Q(operprod[8]) );
  LNQD1BWP \operprod_reg[7]  ( .D(N1926), .EN(N78), .Q(operprod[7]) );
  LNQD1BWP \operprod_reg[6]  ( .D(N1925), .EN(N78), .Q(operprod[6]) );
  LNQD1BWP \operprod_reg[5]  ( .D(N1924), .EN(N78), .Q(operprod[5]) );
  LNQD1BWP \operprod_reg[4]  ( .D(N1923), .EN(N78), .Q(operprod[4]) );
  LNQD1BWP \operprod_reg[3]  ( .D(N1922), .EN(N78), .Q(operprod[3]) );
  LNQD1BWP \operprod_reg[2]  ( .D(N1921), .EN(N78), .Q(operprod[2]) );
  LNQD1BWP \operprod_reg[1]  ( .D(N1920), .EN(N78), .Q(operprod[1]) );
  LNQD1BWP \operprod_reg[0]  ( .D(N1919), .EN(N78), .Q(operprod[0]) );
  LNQD1BWP \temp_exp_reg[6]  ( .D(N1917), .EN(N78), .Q(temp_exp[6]) );
  LNQD1BWP \temp_exp_reg[5]  ( .D(N1916), .EN(N78), .Q(temp_exp[5]) );
  LNQD1BWP \temp_exp_reg[4]  ( .D(N1915), .EN(N78), .Q(temp_exp[4]) );
  LNQD1BWP \temp_exp_reg[3]  ( .D(N1914), .EN(N78), .Q(temp_exp[3]) );
  LNQD1BWP \temp_exp_reg[2]  ( .D(N1913), .EN(N78), .Q(temp_exp[2]) );
  LNQD1BWP \temp_exp_reg[1]  ( .D(N1912), .EN(N78), .Q(temp_exp[1]) );
  LNQD1BWP \temp_exp_reg[0]  ( .D(N1911), .EN(N78), .Q(temp_exp[0]) );
  LHQD1BWP Overflow_reg ( .E(N1942), .D(N78), .Q(Overflow) );
  LHQD1BWP \operprod1_reg[9]  ( .E(n750), .D(N1855), .Q(operprod1[9]) );
  LHQD1BWP \operprod1_reg[8]  ( .E(n750), .D(N1854), .Q(operprod1[8]) );
  LHQD1BWP \operprod1_reg[7]  ( .E(n750), .D(N1853), .Q(operprod1[7]) );
  LHQD1BWP \operprod1_reg[6]  ( .E(n750), .D(N1852), .Q(operprod1[6]) );
  LHQD1BWP \operprod1_reg[5]  ( .E(n750), .D(N1851), .Q(operprod1[5]) );
  LHQD1BWP \operprod1_reg[4]  ( .E(n750), .D(N1850), .Q(operprod1[4]) );
  LHQD1BWP \operprod1_reg[3]  ( .E(n750), .D(N1849), .Q(operprod1[3]) );
  LHQD1BWP \operprod1_reg[2]  ( .E(n750), .D(N1848), .Q(operprod1[2]) );
  LHQD1BWP \operprod1_reg[1]  ( .E(n750), .D(N1847), .Q(operprod1[1]) );
  LHQD1BWP \operprod1_reg[0]  ( .E(n750), .D(N1846), .Q(operprod1[0]) );
  IND2D1BWP \DP_OP_379J1_125_371/U245  ( .A1(B[0]), .B1(A[1]), .ZN(
        \DP_OP_379J1_125_371/n279 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U244  ( .A1(A[1]), .A2(B[0]), .ZN(
        \DP_OP_379J1_125_371/n278 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U243  ( .A1(A[1]), .A2(B[1]), .ZN(
        \DP_OP_379J1_125_371/n277 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U242  ( .A1(A[1]), .A2(B[2]), .ZN(
        \DP_OP_379J1_125_371/n276 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U241  ( .A1(A[1]), .A2(B[3]), .ZN(
        \DP_OP_379J1_125_371/n275 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U240  ( .A1(A[1]), .A2(B[4]), .ZN(
        \DP_OP_379J1_125_371/n274 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U239  ( .A1(A[1]), .A2(B[5]), .ZN(
        \DP_OP_379J1_125_371/n273 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U238  ( .A1(A[1]), .A2(B[6]), .ZN(
        \DP_OP_379J1_125_371/n272 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U237  ( .A1(A[1]), .A2(B[7]), .ZN(
        \DP_OP_379J1_125_371/n271 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U236  ( .A1(A[1]), .A2(B[8]), .ZN(
        \DP_OP_379J1_125_371/n270 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U235  ( .A1(A[1]), .A2(B[9]), .ZN(
        \DP_OP_379J1_125_371/n269 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U234  ( .A1(A[1]), .A2(N93), .ZN(
        \DP_OP_379J1_125_371/n268 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U232  ( .A1(\DP_OP_379J1_125_371/n324 ), 
        .A2(\DP_OP_379J1_125_371/n278 ), .B1(\DP_OP_379J1_125_371/n277 ), .B2(
        n536), .ZN(\DP_OP_379J1_125_371/n208 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U231  ( .A1(\DP_OP_379J1_125_371/n324 ), 
        .A2(\DP_OP_379J1_125_371/n277 ), .B1(\DP_OP_379J1_125_371/n276 ), .B2(
        n536), .ZN(\DP_OP_379J1_125_371/n207 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U230  ( .A1(\DP_OP_379J1_125_371/n324 ), 
        .A2(\DP_OP_379J1_125_371/n276 ), .B1(\DP_OP_379J1_125_371/n275 ), .B2(
        n536), .ZN(\DP_OP_379J1_125_371/n206 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U229  ( .A1(\DP_OP_379J1_125_371/n324 ), 
        .A2(\DP_OP_379J1_125_371/n275 ), .B1(\DP_OP_379J1_125_371/n274 ), .B2(
        n536), .ZN(\DP_OP_379J1_125_371/n205 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U228  ( .A1(\DP_OP_379J1_125_371/n324 ), 
        .A2(\DP_OP_379J1_125_371/n274 ), .B1(\DP_OP_379J1_125_371/n273 ), .B2(
        n536), .ZN(\DP_OP_379J1_125_371/n204 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U227  ( .A1(\DP_OP_379J1_125_371/n324 ), 
        .A2(\DP_OP_379J1_125_371/n273 ), .B1(\DP_OP_379J1_125_371/n272 ), .B2(
        n536), .ZN(\DP_OP_379J1_125_371/n203 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U226  ( .A1(\DP_OP_379J1_125_371/n324 ), 
        .A2(\DP_OP_379J1_125_371/n272 ), .B1(\DP_OP_379J1_125_371/n271 ), .B2(
        n536), .ZN(\DP_OP_379J1_125_371/n202 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U225  ( .A1(\DP_OP_379J1_125_371/n324 ), 
        .A2(\DP_OP_379J1_125_371/n271 ), .B1(\DP_OP_379J1_125_371/n270 ), .B2(
        n536), .ZN(\DP_OP_379J1_125_371/n201 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U224  ( .A1(\DP_OP_379J1_125_371/n324 ), 
        .A2(\DP_OP_379J1_125_371/n270 ), .B1(\DP_OP_379J1_125_371/n269 ), .B2(
        n536), .ZN(\DP_OP_379J1_125_371/n200 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U223  ( .A1(\DP_OP_379J1_125_371/n324 ), 
        .A2(\DP_OP_379J1_125_371/n269 ), .B1(\DP_OP_379J1_125_371/n268 ), .B2(
        n536), .ZN(\DP_OP_379J1_125_371/n199 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U222  ( .A1(\DP_OP_379J1_125_371/n324 ), 
        .A2(\DP_OP_379J1_125_371/n268 ), .B1(n537), .B2(n536), .ZN(
        \DP_OP_379J1_125_371/n198 ) );
  AO21D1BWP \DP_OP_379J1_125_371/U221  ( .A1(\DP_OP_379J1_125_371/n324 ), .A2(
        n536), .B(n537), .Z(\DP_OP_379J1_125_371/n197 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U220  ( .A1(\DP_OP_379J1_125_371/n324 ), 
        .A2(n537), .B1(\DP_OP_379J1_125_371/n279 ), .B2(n536), .ZN(
        \DP_OP_379J1_125_371/n136 ) );
  IND2D1BWP \DP_OP_379J1_125_371/U219  ( .A1(B[0]), .B1(A[3]), .ZN(
        \DP_OP_379J1_125_371/n267 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U218  ( .A1(A[3]), .A2(B[0]), .ZN(
        \DP_OP_379J1_125_371/n266 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U217  ( .A1(A[3]), .A2(B[1]), .ZN(
        \DP_OP_379J1_125_371/n265 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U216  ( .A1(A[3]), .A2(B[2]), .ZN(
        \DP_OP_379J1_125_371/n264 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U215  ( .A1(A[3]), .A2(B[3]), .ZN(
        \DP_OP_379J1_125_371/n263 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U214  ( .A1(A[3]), .A2(B[4]), .ZN(
        \DP_OP_379J1_125_371/n262 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U213  ( .A1(A[3]), .A2(B[5]), .ZN(
        \DP_OP_379J1_125_371/n261 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U212  ( .A1(A[3]), .A2(B[6]), .ZN(
        \DP_OP_379J1_125_371/n260 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U211  ( .A1(A[3]), .A2(B[7]), .ZN(
        \DP_OP_379J1_125_371/n259 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U210  ( .A1(A[3]), .A2(B[8]), .ZN(
        \DP_OP_379J1_125_371/n258 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U209  ( .A1(A[3]), .A2(B[9]), .ZN(
        \DP_OP_379J1_125_371/n257 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U208  ( .A1(A[3]), .A2(N93), .ZN(
        \DP_OP_379J1_125_371/n256 ) );
  INR2D1BWP \DP_OP_379J1_125_371/U207  ( .A1(B[0]), .B1(
        \DP_OP_379J1_125_371/n329 ), .ZN(\DP_OP_379J1_125_371/n196 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U206  ( .A1(\DP_OP_379J1_125_371/n323 ), 
        .A2(\DP_OP_379J1_125_371/n266 ), .B1(\DP_OP_379J1_125_371/n329 ), .B2(
        \DP_OP_379J1_125_371/n265 ), .ZN(\DP_OP_379J1_125_371/n195 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U205  ( .A1(\DP_OP_379J1_125_371/n323 ), 
        .A2(\DP_OP_379J1_125_371/n265 ), .B1(\DP_OP_379J1_125_371/n329 ), .B2(
        \DP_OP_379J1_125_371/n264 ), .ZN(\DP_OP_379J1_125_371/n194 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U204  ( .A1(\DP_OP_379J1_125_371/n323 ), 
        .A2(\DP_OP_379J1_125_371/n264 ), .B1(\DP_OP_379J1_125_371/n329 ), .B2(
        \DP_OP_379J1_125_371/n263 ), .ZN(\DP_OP_379J1_125_371/n193 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U203  ( .A1(\DP_OP_379J1_125_371/n323 ), 
        .A2(\DP_OP_379J1_125_371/n263 ), .B1(\DP_OP_379J1_125_371/n329 ), .B2(
        \DP_OP_379J1_125_371/n262 ), .ZN(\DP_OP_379J1_125_371/n192 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U202  ( .A1(\DP_OP_379J1_125_371/n323 ), 
        .A2(\DP_OP_379J1_125_371/n262 ), .B1(\DP_OP_379J1_125_371/n329 ), .B2(
        \DP_OP_379J1_125_371/n261 ), .ZN(\DP_OP_379J1_125_371/n191 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U201  ( .A1(\DP_OP_379J1_125_371/n323 ), 
        .A2(\DP_OP_379J1_125_371/n261 ), .B1(\DP_OP_379J1_125_371/n329 ), .B2(
        \DP_OP_379J1_125_371/n260 ), .ZN(\DP_OP_379J1_125_371/n190 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U200  ( .A1(\DP_OP_379J1_125_371/n323 ), 
        .A2(\DP_OP_379J1_125_371/n260 ), .B1(\DP_OP_379J1_125_371/n329 ), .B2(
        \DP_OP_379J1_125_371/n259 ), .ZN(\DP_OP_379J1_125_371/n189 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U199  ( .A1(\DP_OP_379J1_125_371/n323 ), 
        .A2(\DP_OP_379J1_125_371/n259 ), .B1(\DP_OP_379J1_125_371/n329 ), .B2(
        \DP_OP_379J1_125_371/n258 ), .ZN(\DP_OP_379J1_125_371/n188 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U198  ( .A1(\DP_OP_379J1_125_371/n323 ), 
        .A2(\DP_OP_379J1_125_371/n258 ), .B1(\DP_OP_379J1_125_371/n329 ), .B2(
        \DP_OP_379J1_125_371/n257 ), .ZN(\DP_OP_379J1_125_371/n187 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U197  ( .A1(\DP_OP_379J1_125_371/n323 ), 
        .A2(\DP_OP_379J1_125_371/n257 ), .B1(\DP_OP_379J1_125_371/n329 ), .B2(
        \DP_OP_379J1_125_371/n256 ), .ZN(\DP_OP_379J1_125_371/n186 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U196  ( .A1(\DP_OP_379J1_125_371/n323 ), 
        .A2(\DP_OP_379J1_125_371/n256 ), .B1(\DP_OP_379J1_125_371/n329 ), .B2(
        n538), .ZN(\DP_OP_379J1_125_371/n185 ) );
  AO21D1BWP \DP_OP_379J1_125_371/U195  ( .A1(\DP_OP_379J1_125_371/n323 ), .A2(
        \DP_OP_379J1_125_371/n329 ), .B(n538), .Z(\DP_OP_379J1_125_371/n184 )
         );
  OAI22D1BWP \DP_OP_379J1_125_371/U194  ( .A1(\DP_OP_379J1_125_371/n323 ), 
        .A2(n538), .B1(\DP_OP_379J1_125_371/n329 ), .B2(
        \DP_OP_379J1_125_371/n267 ), .ZN(\DP_OP_379J1_125_371/n135 ) );
  IND2D1BWP \DP_OP_379J1_125_371/U193  ( .A1(B[0]), .B1(A[5]), .ZN(
        \DP_OP_379J1_125_371/n255 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U192  ( .A1(A[5]), .A2(B[0]), .ZN(
        \DP_OP_379J1_125_371/n254 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U191  ( .A1(A[5]), .A2(B[1]), .ZN(
        \DP_OP_379J1_125_371/n253 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U190  ( .A1(A[5]), .A2(B[2]), .ZN(
        \DP_OP_379J1_125_371/n252 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U189  ( .A1(A[5]), .A2(B[3]), .ZN(
        \DP_OP_379J1_125_371/n251 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U188  ( .A1(A[5]), .A2(B[4]), .ZN(
        \DP_OP_379J1_125_371/n250 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U187  ( .A1(A[5]), .A2(B[5]), .ZN(
        \DP_OP_379J1_125_371/n249 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U186  ( .A1(A[5]), .A2(B[6]), .ZN(
        \DP_OP_379J1_125_371/n248 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U185  ( .A1(A[5]), .A2(B[7]), .ZN(
        \DP_OP_379J1_125_371/n247 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U184  ( .A1(A[5]), .A2(B[8]), .ZN(
        \DP_OP_379J1_125_371/n246 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U183  ( .A1(A[5]), .A2(B[9]), .ZN(
        \DP_OP_379J1_125_371/n245 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U182  ( .A1(A[5]), .A2(N93), .ZN(
        \DP_OP_379J1_125_371/n244 ) );
  INR2D1BWP \DP_OP_379J1_125_371/U181  ( .A1(B[0]), .B1(
        \DP_OP_379J1_125_371/n328 ), .ZN(\DP_OP_379J1_125_371/n183 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U180  ( .A1(\DP_OP_379J1_125_371/n322 ), 
        .A2(\DP_OP_379J1_125_371/n254 ), .B1(\DP_OP_379J1_125_371/n328 ), .B2(
        \DP_OP_379J1_125_371/n253 ), .ZN(\DP_OP_379J1_125_371/n182 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U179  ( .A1(\DP_OP_379J1_125_371/n322 ), 
        .A2(\DP_OP_379J1_125_371/n253 ), .B1(\DP_OP_379J1_125_371/n328 ), .B2(
        \DP_OP_379J1_125_371/n252 ), .ZN(\DP_OP_379J1_125_371/n181 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U178  ( .A1(\DP_OP_379J1_125_371/n322 ), 
        .A2(\DP_OP_379J1_125_371/n252 ), .B1(\DP_OP_379J1_125_371/n328 ), .B2(
        \DP_OP_379J1_125_371/n251 ), .ZN(\DP_OP_379J1_125_371/n180 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U177  ( .A1(\DP_OP_379J1_125_371/n322 ), 
        .A2(\DP_OP_379J1_125_371/n251 ), .B1(\DP_OP_379J1_125_371/n328 ), .B2(
        \DP_OP_379J1_125_371/n250 ), .ZN(\DP_OP_379J1_125_371/n179 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U176  ( .A1(\DP_OP_379J1_125_371/n322 ), 
        .A2(\DP_OP_379J1_125_371/n250 ), .B1(\DP_OP_379J1_125_371/n328 ), .B2(
        \DP_OP_379J1_125_371/n249 ), .ZN(\DP_OP_379J1_125_371/n178 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U175  ( .A1(\DP_OP_379J1_125_371/n322 ), 
        .A2(\DP_OP_379J1_125_371/n249 ), .B1(\DP_OP_379J1_125_371/n328 ), .B2(
        \DP_OP_379J1_125_371/n248 ), .ZN(\DP_OP_379J1_125_371/n177 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U174  ( .A1(\DP_OP_379J1_125_371/n322 ), 
        .A2(\DP_OP_379J1_125_371/n248 ), .B1(\DP_OP_379J1_125_371/n328 ), .B2(
        \DP_OP_379J1_125_371/n247 ), .ZN(\DP_OP_379J1_125_371/n176 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U173  ( .A1(\DP_OP_379J1_125_371/n322 ), 
        .A2(\DP_OP_379J1_125_371/n247 ), .B1(\DP_OP_379J1_125_371/n328 ), .B2(
        \DP_OP_379J1_125_371/n246 ), .ZN(\DP_OP_379J1_125_371/n175 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U172  ( .A1(\DP_OP_379J1_125_371/n322 ), 
        .A2(\DP_OP_379J1_125_371/n246 ), .B1(\DP_OP_379J1_125_371/n328 ), .B2(
        \DP_OP_379J1_125_371/n245 ), .ZN(\DP_OP_379J1_125_371/n174 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U171  ( .A1(\DP_OP_379J1_125_371/n322 ), 
        .A2(\DP_OP_379J1_125_371/n245 ), .B1(\DP_OP_379J1_125_371/n328 ), .B2(
        \DP_OP_379J1_125_371/n244 ), .ZN(\DP_OP_379J1_125_371/n173 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U170  ( .A1(\DP_OP_379J1_125_371/n322 ), 
        .A2(\DP_OP_379J1_125_371/n244 ), .B1(\DP_OP_379J1_125_371/n328 ), .B2(
        n539), .ZN(\DP_OP_379J1_125_371/n172 ) );
  AO21D1BWP \DP_OP_379J1_125_371/U169  ( .A1(\DP_OP_379J1_125_371/n322 ), .A2(
        \DP_OP_379J1_125_371/n328 ), .B(n539), .Z(\DP_OP_379J1_125_371/n171 )
         );
  OAI22D1BWP \DP_OP_379J1_125_371/U168  ( .A1(\DP_OP_379J1_125_371/n322 ), 
        .A2(n539), .B1(\DP_OP_379J1_125_371/n328 ), .B2(
        \DP_OP_379J1_125_371/n255 ), .ZN(\DP_OP_379J1_125_371/n134 ) );
  IND2D1BWP \DP_OP_379J1_125_371/U167  ( .A1(B[0]), .B1(A[7]), .ZN(
        \DP_OP_379J1_125_371/n243 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U166  ( .A1(A[7]), .A2(B[0]), .ZN(
        \DP_OP_379J1_125_371/n242 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U165  ( .A1(A[7]), .A2(B[1]), .ZN(
        \DP_OP_379J1_125_371/n241 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U164  ( .A1(A[7]), .A2(B[2]), .ZN(
        \DP_OP_379J1_125_371/n240 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U163  ( .A1(A[7]), .A2(B[3]), .ZN(
        \DP_OP_379J1_125_371/n239 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U162  ( .A1(A[7]), .A2(B[4]), .ZN(
        \DP_OP_379J1_125_371/n238 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U161  ( .A1(A[7]), .A2(B[5]), .ZN(
        \DP_OP_379J1_125_371/n237 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U160  ( .A1(A[7]), .A2(B[6]), .ZN(
        \DP_OP_379J1_125_371/n236 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U159  ( .A1(A[7]), .A2(B[7]), .ZN(
        \DP_OP_379J1_125_371/n235 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U158  ( .A1(A[7]), .A2(B[8]), .ZN(
        \DP_OP_379J1_125_371/n234 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U157  ( .A1(A[7]), .A2(B[9]), .ZN(
        \DP_OP_379J1_125_371/n233 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U156  ( .A1(A[7]), .A2(N93), .ZN(
        \DP_OP_379J1_125_371/n232 ) );
  INR2D1BWP \DP_OP_379J1_125_371/U155  ( .A1(B[0]), .B1(
        \DP_OP_379J1_125_371/n327 ), .ZN(\DP_OP_379J1_125_371/n170 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U154  ( .A1(\DP_OP_379J1_125_371/n321 ), 
        .A2(\DP_OP_379J1_125_371/n242 ), .B1(\DP_OP_379J1_125_371/n327 ), .B2(
        \DP_OP_379J1_125_371/n241 ), .ZN(\DP_OP_379J1_125_371/n169 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U153  ( .A1(\DP_OP_379J1_125_371/n321 ), 
        .A2(\DP_OP_379J1_125_371/n241 ), .B1(\DP_OP_379J1_125_371/n327 ), .B2(
        \DP_OP_379J1_125_371/n240 ), .ZN(\DP_OP_379J1_125_371/n168 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U152  ( .A1(\DP_OP_379J1_125_371/n321 ), 
        .A2(\DP_OP_379J1_125_371/n240 ), .B1(\DP_OP_379J1_125_371/n327 ), .B2(
        \DP_OP_379J1_125_371/n239 ), .ZN(\DP_OP_379J1_125_371/n167 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U151  ( .A1(\DP_OP_379J1_125_371/n321 ), 
        .A2(\DP_OP_379J1_125_371/n239 ), .B1(\DP_OP_379J1_125_371/n327 ), .B2(
        \DP_OP_379J1_125_371/n238 ), .ZN(\DP_OP_379J1_125_371/n166 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U150  ( .A1(\DP_OP_379J1_125_371/n321 ), 
        .A2(\DP_OP_379J1_125_371/n238 ), .B1(\DP_OP_379J1_125_371/n327 ), .B2(
        \DP_OP_379J1_125_371/n237 ), .ZN(\DP_OP_379J1_125_371/n165 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U149  ( .A1(\DP_OP_379J1_125_371/n321 ), 
        .A2(\DP_OP_379J1_125_371/n237 ), .B1(\DP_OP_379J1_125_371/n327 ), .B2(
        \DP_OP_379J1_125_371/n236 ), .ZN(\DP_OP_379J1_125_371/n164 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U148  ( .A1(\DP_OP_379J1_125_371/n321 ), 
        .A2(\DP_OP_379J1_125_371/n236 ), .B1(\DP_OP_379J1_125_371/n327 ), .B2(
        \DP_OP_379J1_125_371/n235 ), .ZN(\DP_OP_379J1_125_371/n163 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U147  ( .A1(\DP_OP_379J1_125_371/n321 ), 
        .A2(\DP_OP_379J1_125_371/n235 ), .B1(\DP_OP_379J1_125_371/n327 ), .B2(
        \DP_OP_379J1_125_371/n234 ), .ZN(\DP_OP_379J1_125_371/n162 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U146  ( .A1(\DP_OP_379J1_125_371/n321 ), 
        .A2(\DP_OP_379J1_125_371/n234 ), .B1(\DP_OP_379J1_125_371/n327 ), .B2(
        \DP_OP_379J1_125_371/n233 ), .ZN(\DP_OP_379J1_125_371/n161 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U145  ( .A1(\DP_OP_379J1_125_371/n321 ), 
        .A2(\DP_OP_379J1_125_371/n233 ), .B1(\DP_OP_379J1_125_371/n327 ), .B2(
        \DP_OP_379J1_125_371/n232 ), .ZN(\DP_OP_379J1_125_371/n160 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U144  ( .A1(\DP_OP_379J1_125_371/n321 ), 
        .A2(\DP_OP_379J1_125_371/n232 ), .B1(\DP_OP_379J1_125_371/n327 ), .B2(
        n540), .ZN(\DP_OP_379J1_125_371/n159 ) );
  AO21D1BWP \DP_OP_379J1_125_371/U143  ( .A1(\DP_OP_379J1_125_371/n321 ), .A2(
        \DP_OP_379J1_125_371/n327 ), .B(n540), .Z(\DP_OP_379J1_125_371/n158 )
         );
  OAI22D1BWP \DP_OP_379J1_125_371/U142  ( .A1(\DP_OP_379J1_125_371/n321 ), 
        .A2(n540), .B1(\DP_OP_379J1_125_371/n327 ), .B2(
        \DP_OP_379J1_125_371/n243 ), .ZN(\DP_OP_379J1_125_371/n133 ) );
  IND2D1BWP \DP_OP_379J1_125_371/U141  ( .A1(B[0]), .B1(A[9]), .ZN(
        \DP_OP_379J1_125_371/n231 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U140  ( .A1(A[9]), .A2(B[0]), .ZN(
        \DP_OP_379J1_125_371/n230 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U139  ( .A1(A[9]), .A2(B[1]), .ZN(
        \DP_OP_379J1_125_371/n229 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U138  ( .A1(A[9]), .A2(B[2]), .ZN(
        \DP_OP_379J1_125_371/n228 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U137  ( .A1(A[9]), .A2(B[3]), .ZN(
        \DP_OP_379J1_125_371/n227 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U136  ( .A1(A[9]), .A2(B[4]), .ZN(
        \DP_OP_379J1_125_371/n226 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U135  ( .A1(A[9]), .A2(B[5]), .ZN(
        \DP_OP_379J1_125_371/n225 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U134  ( .A1(A[9]), .A2(B[6]), .ZN(
        \DP_OP_379J1_125_371/n224 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U133  ( .A1(A[9]), .A2(B[7]), .ZN(
        \DP_OP_379J1_125_371/n223 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U132  ( .A1(A[9]), .A2(B[8]), .ZN(
        \DP_OP_379J1_125_371/n222 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U131  ( .A1(A[9]), .A2(B[9]), .ZN(
        \DP_OP_379J1_125_371/n221 ) );
  XNR2D1BWP \DP_OP_379J1_125_371/U130  ( .A1(A[9]), .A2(N93), .ZN(
        \DP_OP_379J1_125_371/n220 ) );
  INR2D1BWP \DP_OP_379J1_125_371/U129  ( .A1(B[0]), .B1(
        \DP_OP_379J1_125_371/n326 ), .ZN(\DP_OP_379J1_125_371/n157 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U128  ( .A1(\DP_OP_379J1_125_371/n320 ), 
        .A2(\DP_OP_379J1_125_371/n230 ), .B1(\DP_OP_379J1_125_371/n326 ), .B2(
        \DP_OP_379J1_125_371/n229 ), .ZN(\DP_OP_379J1_125_371/n156 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U127  ( .A1(\DP_OP_379J1_125_371/n320 ), 
        .A2(\DP_OP_379J1_125_371/n229 ), .B1(\DP_OP_379J1_125_371/n326 ), .B2(
        \DP_OP_379J1_125_371/n228 ), .ZN(\DP_OP_379J1_125_371/n155 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U126  ( .A1(\DP_OP_379J1_125_371/n320 ), 
        .A2(\DP_OP_379J1_125_371/n228 ), .B1(\DP_OP_379J1_125_371/n326 ), .B2(
        \DP_OP_379J1_125_371/n227 ), .ZN(\DP_OP_379J1_125_371/n154 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U125  ( .A1(\DP_OP_379J1_125_371/n320 ), 
        .A2(\DP_OP_379J1_125_371/n227 ), .B1(\DP_OP_379J1_125_371/n326 ), .B2(
        \DP_OP_379J1_125_371/n226 ), .ZN(\DP_OP_379J1_125_371/n153 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U124  ( .A1(\DP_OP_379J1_125_371/n320 ), 
        .A2(\DP_OP_379J1_125_371/n226 ), .B1(\DP_OP_379J1_125_371/n326 ), .B2(
        \DP_OP_379J1_125_371/n225 ), .ZN(\DP_OP_379J1_125_371/n152 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U123  ( .A1(\DP_OP_379J1_125_371/n320 ), 
        .A2(\DP_OP_379J1_125_371/n225 ), .B1(\DP_OP_379J1_125_371/n326 ), .B2(
        \DP_OP_379J1_125_371/n224 ), .ZN(\DP_OP_379J1_125_371/n151 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U122  ( .A1(\DP_OP_379J1_125_371/n320 ), 
        .A2(\DP_OP_379J1_125_371/n224 ), .B1(\DP_OP_379J1_125_371/n326 ), .B2(
        \DP_OP_379J1_125_371/n223 ), .ZN(\DP_OP_379J1_125_371/n150 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U121  ( .A1(\DP_OP_379J1_125_371/n320 ), 
        .A2(\DP_OP_379J1_125_371/n223 ), .B1(\DP_OP_379J1_125_371/n326 ), .B2(
        \DP_OP_379J1_125_371/n222 ), .ZN(\DP_OP_379J1_125_371/n149 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U120  ( .A1(\DP_OP_379J1_125_371/n320 ), 
        .A2(\DP_OP_379J1_125_371/n222 ), .B1(\DP_OP_379J1_125_371/n326 ), .B2(
        \DP_OP_379J1_125_371/n221 ), .ZN(\DP_OP_379J1_125_371/n148 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U119  ( .A1(\DP_OP_379J1_125_371/n320 ), 
        .A2(\DP_OP_379J1_125_371/n221 ), .B1(\DP_OP_379J1_125_371/n326 ), .B2(
        \DP_OP_379J1_125_371/n220 ), .ZN(\DP_OP_379J1_125_371/n147 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U118  ( .A1(\DP_OP_379J1_125_371/n320 ), 
        .A2(\DP_OP_379J1_125_371/n220 ), .B1(\DP_OP_379J1_125_371/n326 ), .B2(
        n541), .ZN(\DP_OP_379J1_125_371/n146 ) );
  AO21D1BWP \DP_OP_379J1_125_371/U117  ( .A1(\DP_OP_379J1_125_371/n320 ), .A2(
        \DP_OP_379J1_125_371/n326 ), .B(n541), .Z(\DP_OP_379J1_125_371/n145 )
         );
  OAI22D1BWP \DP_OP_379J1_125_371/U116  ( .A1(\DP_OP_379J1_125_371/n320 ), 
        .A2(n541), .B1(\DP_OP_379J1_125_371/n326 ), .B2(
        \DP_OP_379J1_125_371/n231 ), .ZN(\DP_OP_379J1_125_371/n132 ) );
  INR2D1BWP \DP_OP_379J1_125_371/U104  ( .A1(B[0]), .B1(
        \DP_OP_379J1_125_371/n325 ), .ZN(\DP_OP_379J1_125_371/n144 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U103  ( .A1(\DP_OP_379J1_125_371/n319 ), 
        .A2(n525), .B1(\DP_OP_379J1_125_371/n325 ), .B2(n526), .ZN(
        \DP_OP_379J1_125_371/n143 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U102  ( .A1(\DP_OP_379J1_125_371/n319 ), 
        .A2(n526), .B1(\DP_OP_379J1_125_371/n325 ), .B2(n527), .ZN(
        \DP_OP_379J1_125_371/n83 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U101  ( .A1(\DP_OP_379J1_125_371/n319 ), 
        .A2(n527), .B1(\DP_OP_379J1_125_371/n325 ), .B2(n528), .ZN(
        \DP_OP_379J1_125_371/n142 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U100  ( .A1(\DP_OP_379J1_125_371/n319 ), 
        .A2(n528), .B1(\DP_OP_379J1_125_371/n325 ), .B2(n529), .ZN(
        \DP_OP_379J1_125_371/n141 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U99  ( .A1(\DP_OP_379J1_125_371/n319 ), .A2(
        n529), .B1(\DP_OP_379J1_125_371/n325 ), .B2(n530), .ZN(
        \DP_OP_379J1_125_371/n69 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U98  ( .A1(\DP_OP_379J1_125_371/n319 ), .A2(
        n530), .B1(\DP_OP_379J1_125_371/n325 ), .B2(n531), .ZN(
        \DP_OP_379J1_125_371/n140 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U97  ( .A1(\DP_OP_379J1_125_371/n319 ), .A2(
        n531), .B1(\DP_OP_379J1_125_371/n325 ), .B2(n532), .ZN(
        \DP_OP_379J1_125_371/n57 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U96  ( .A1(\DP_OP_379J1_125_371/n319 ), .A2(
        n532), .B1(\DP_OP_379J1_125_371/n325 ), .B2(n533), .ZN(
        \DP_OP_379J1_125_371/n139 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U94  ( .A1(\DP_OP_379J1_125_371/n319 ), .A2(
        n534), .B1(\DP_OP_379J1_125_371/n325 ), .B2(n535), .ZN(
        \DP_OP_379J1_125_371/n138 ) );
  FA1D0BWP \DP_OP_379J1_125_371/U91  ( .A(\DP_OP_379J1_125_371/n205 ), .B(
        \DP_OP_379J1_125_371/n183 ), .CI(\DP_OP_379J1_125_371/n194 ), .CO(
        \DP_OP_379J1_125_371/n128 ), .S(\DP_OP_379J1_125_371/n129 ) );
  FA1D0BWP \DP_OP_379J1_125_371/U89  ( .A(\DP_OP_379J1_125_371/n193 ), .B(
        \DP_OP_379J1_125_371/n204 ), .CI(\DP_OP_379J1_125_371/n127 ), .CO(
        \DP_OP_379J1_125_371/n124 ), .S(\DP_OP_379J1_125_371/n125 ) );
  CMPE42D1BWP \DP_OP_379J1_125_371/U88  ( .A(\DP_OP_379J1_125_371/n203 ), .B(
        \DP_OP_379J1_125_371/n170 ), .C(\DP_OP_379J1_125_371/n181 ), .CIX(
        \DP_OP_379J1_125_371/n126 ), .D(\DP_OP_379J1_125_371/n192 ), .CO(
        \DP_OP_379J1_125_371/n122 ), .COX(\DP_OP_379J1_125_371/n121 ), .S(
        \DP_OP_379J1_125_371/n123 ) );
  CMPE42D1BWP \DP_OP_379J1_125_371/U86  ( .A(\DP_OP_379J1_125_371/n180 ), .B(
        \DP_OP_379J1_125_371/n202 ), .C(\DP_OP_379J1_125_371/n191 ), .CIX(
        \DP_OP_379J1_125_371/n121 ), .D(\DP_OP_379J1_125_371/n120 ), .CO(
        \DP_OP_379J1_125_371/n117 ), .COX(\DP_OP_379J1_125_371/n116 ), .S(
        \DP_OP_379J1_125_371/n118 ) );
  FA1D0BWP \DP_OP_379J1_125_371/U85  ( .A(\DP_OP_379J1_125_371/n179 ), .B(
        \DP_OP_379J1_125_371/n157 ), .CI(\DP_OP_379J1_125_371/n168 ), .CO(
        \DP_OP_379J1_125_371/n114 ), .S(\DP_OP_379J1_125_371/n115 ) );
  CMPE42D1BWP \DP_OP_379J1_125_371/U84  ( .A(\DP_OP_379J1_125_371/n190 ), .B(
        \DP_OP_379J1_125_371/n201 ), .C(\DP_OP_379J1_125_371/n119 ), .CIX(
        \DP_OP_379J1_125_371/n115 ), .D(\DP_OP_379J1_125_371/n116 ), .CO(
        \DP_OP_379J1_125_371/n112 ), .COX(\DP_OP_379J1_125_371/n111 ), .S(
        \DP_OP_379J1_125_371/n113 ) );
  FA1D0BWP \DP_OP_379J1_125_371/U82  ( .A(\DP_OP_379J1_125_371/n167 ), .B(
        \DP_OP_379J1_125_371/n178 ), .CI(\DP_OP_379J1_125_371/n189 ), .CO(
        \DP_OP_379J1_125_371/n107 ), .S(\DP_OP_379J1_125_371/n108 ) );
  CMPE42D1BWP \DP_OP_379J1_125_371/U81  ( .A(\DP_OP_379J1_125_371/n110 ), .B(
        \DP_OP_379J1_125_371/n200 ), .C(\DP_OP_379J1_125_371/n114 ), .CIX(
        \DP_OP_379J1_125_371/n111 ), .D(\DP_OP_379J1_125_371/n108 ), .CO(
        \DP_OP_379J1_125_371/n105 ), .COX(\DP_OP_379J1_125_371/n104 ), .S(
        \DP_OP_379J1_125_371/n106 ) );
  CMPE42D1BWP \DP_OP_379J1_125_371/U80  ( .A(\DP_OP_379J1_125_371/n166 ), .B(
        \DP_OP_379J1_125_371/n144 ), .C(\DP_OP_379J1_125_371/n155 ), .CIX(
        \DP_OP_379J1_125_371/n107 ), .D(\DP_OP_379J1_125_371/n177 ), .CO(
        \DP_OP_379J1_125_371/n102 ), .COX(\DP_OP_379J1_125_371/n101 ), .S(
        \DP_OP_379J1_125_371/n103 ) );
  CMPE42D1BWP \DP_OP_379J1_125_371/U79  ( .A(\DP_OP_379J1_125_371/n188 ), .B(
        \DP_OP_379J1_125_371/n199 ), .C(\DP_OP_379J1_125_371/n109 ), .CIX(
        \DP_OP_379J1_125_371/n103 ), .D(\DP_OP_379J1_125_371/n104 ), .CO(
        \DP_OP_379J1_125_371/n99 ), .COX(\DP_OP_379J1_125_371/n98 ), .S(
        \DP_OP_379J1_125_371/n100 ) );
  CMPE42D1BWP \DP_OP_379J1_125_371/U78  ( .A(\DP_OP_379J1_125_371/n154 ), .B(
        \DP_OP_379J1_125_371/n143 ), .C(\DP_OP_379J1_125_371/n165 ), .CIX(
        \DP_OP_379J1_125_371/n98 ), .D(\DP_OP_379J1_125_371/n176 ), .CO(
        \DP_OP_379J1_125_371/n96 ), .COX(\DP_OP_379J1_125_371/n95 ), .S(
        \DP_OP_379J1_125_371/n97 ) );
  CMPE42D1BWP \DP_OP_379J1_125_371/U77  ( .A(\DP_OP_379J1_125_371/n187 ), .B(
        \DP_OP_379J1_125_371/n198 ), .C(\DP_OP_379J1_125_371/n101 ), .CIX(
        \DP_OP_379J1_125_371/n102 ), .D(\DP_OP_379J1_125_371/n97 ), .CO(
        \DP_OP_379J1_125_371/n93 ), .COX(\DP_OP_379J1_125_371/n92 ), .S(
        \DP_OP_379J1_125_371/n94 ) );
  CMPE42D1BWP \DP_OP_379J1_125_371/U75  ( .A(\DP_OP_379J1_125_371/n153 ), .B(
        \DP_OP_379J1_125_371/n175 ), .C(\DP_OP_379J1_125_371/n197 ), .CIX(
        \DP_OP_379J1_125_371/n95 ), .D(n542), .CO(\DP_OP_379J1_125_371/n89 ), 
        .COX(\DP_OP_379J1_125_371/n88 ), .S(\DP_OP_379J1_125_371/n90 ) );
  CMPE42D1BWP \DP_OP_379J1_125_371/U74  ( .A(\DP_OP_379J1_125_371/n164 ), .B(
        \DP_OP_379J1_125_371/n186 ), .C(\DP_OP_379J1_125_371/n92 ), .CIX(
        \DP_OP_379J1_125_371/n96 ), .D(\DP_OP_379J1_125_371/n90 ), .CO(
        \DP_OP_379J1_125_371/n86 ), .COX(\DP_OP_379J1_125_371/n85 ), .S(
        \DP_OP_379J1_125_371/n87 ) );
  CMPE42D1BWP \DP_OP_379J1_125_371/U72  ( .A(\DP_OP_379J1_125_371/n185 ), .B(
        \DP_OP_379J1_125_371/n142 ), .C(\DP_OP_379J1_125_371/n152 ), .CIX(
        \DP_OP_379J1_125_371/n88 ), .D(n542), .CO(\DP_OP_379J1_125_371/n81 ), 
        .COX(\DP_OP_379J1_125_371/n80 ), .S(\DP_OP_379J1_125_371/n82 ) );
  CMPE42D1BWP \DP_OP_379J1_125_371/U71  ( .A(\DP_OP_379J1_125_371/n163 ), .B(
        \DP_OP_379J1_125_371/n174 ), .C(\DP_OP_379J1_125_371/n82 ), .CIX(
        \DP_OP_379J1_125_371/n89 ), .D(\DP_OP_379J1_125_371/n85 ), .CO(
        \DP_OP_379J1_125_371/n78 ), .COX(\DP_OP_379J1_125_371/n77 ), .S(
        \DP_OP_379J1_125_371/n79 ) );
  CMPE42D1BWP \DP_OP_379J1_125_371/U70  ( .A(\DP_OP_379J1_125_371/n173 ), .B(
        \DP_OP_379J1_125_371/n83 ), .C(\DP_OP_379J1_125_371/n162 ), .CIX(
        \DP_OP_379J1_125_371/n80 ), .D(\DP_OP_379J1_125_371/n184 ), .CO(
        \DP_OP_379J1_125_371/n75 ), .COX(\DP_OP_379J1_125_371/n74 ), .S(
        \DP_OP_379J1_125_371/n76 ) );
  CMPE42D1BWP \DP_OP_379J1_125_371/U69  ( .A(\DP_OP_379J1_125_371/n151 ), .B(
        \DP_OP_379J1_125_371/n141 ), .C(\DP_OP_379J1_125_371/n76 ), .CIX(
        \DP_OP_379J1_125_371/n77 ), .D(\DP_OP_379J1_125_371/n81 ), .CO(
        \DP_OP_379J1_125_371/n72 ), .COX(\DP_OP_379J1_125_371/n71 ), .S(
        \DP_OP_379J1_125_371/n73 ) );
  FA1D0BWP \DP_OP_379J1_125_371/U67  ( .A(\DP_OP_379J1_125_371/n161 ), .B(
        \DP_OP_379J1_125_371/n150 ), .CI(n543), .CO(\DP_OP_379J1_125_371/n67 ), 
        .S(\DP_OP_379J1_125_371/n68 ) );
  CMPE42D1BWP \DP_OP_379J1_125_371/U66  ( .A(\DP_OP_379J1_125_371/n74 ), .B(
        \DP_OP_379J1_125_371/n172 ), .C(\DP_OP_379J1_125_371/n68 ), .CIX(
        \DP_OP_379J1_125_371/n71 ), .D(\DP_OP_379J1_125_371/n75 ), .CO(
        \DP_OP_379J1_125_371/n65 ), .COX(\DP_OP_379J1_125_371/n64 ), .S(
        \DP_OP_379J1_125_371/n66 ) );
  FA1D0BWP \DP_OP_379J1_125_371/U65  ( .A(\DP_OP_379J1_125_371/n149 ), .B(
        \DP_OP_379J1_125_371/n69 ), .CI(\DP_OP_379J1_125_371/n171 ), .CO(
        \DP_OP_379J1_125_371/n62 ), .S(\DP_OP_379J1_125_371/n63 ) );
  CMPE42D1BWP \DP_OP_379J1_125_371/U64  ( .A(\DP_OP_379J1_125_371/n160 ), .B(
        \DP_OP_379J1_125_371/n140 ), .C(\DP_OP_379J1_125_371/n67 ), .CIX(
        \DP_OP_379J1_125_371/n64 ), .D(\DP_OP_379J1_125_371/n63 ), .CO(
        \DP_OP_379J1_125_371/n60 ), .COX(\DP_OP_379J1_125_371/n59 ), .S(
        \DP_OP_379J1_125_371/n61 ) );
  CMPE42D1BWP \DP_OP_379J1_125_371/U62  ( .A(\DP_OP_379J1_125_371/n148 ), .B(
        \DP_OP_379J1_125_371/n159 ), .C(n544), .CIX(\DP_OP_379J1_125_371/n59 ), 
        .D(\DP_OP_379J1_125_371/n62 ), .CO(\DP_OP_379J1_125_371/n55 ), .COX(
        \DP_OP_379J1_125_371/n54 ), .S(\DP_OP_379J1_125_371/n56 ) );
  CMPE42D1BWP \DP_OP_379J1_125_371/U61  ( .A(\DP_OP_379J1_125_371/n139 ), .B(
        \DP_OP_379J1_125_371/n57 ), .C(\DP_OP_379J1_125_371/n147 ), .CIX(
        \DP_OP_379J1_125_371/n54 ), .D(\DP_OP_379J1_125_371/n158 ), .CO(
        \DP_OP_379J1_125_371/n52 ), .COX(\DP_OP_379J1_125_371/n51 ), .S(
        \DP_OP_379J1_125_371/n53 ) );
  FA1D0BWP \DP_OP_379J1_125_371/U59  ( .A(n545), .B(\DP_OP_379J1_125_371/n146 ), .CI(\DP_OP_379J1_125_371/n51 ), .CO(\DP_OP_379J1_125_371/n47 ), .S(
        \DP_OP_379J1_125_371/n48 ) );
  FA1D0BWP \DP_OP_379J1_125_371/U55  ( .A(\DP_OP_379J1_125_371/n207 ), .B(
        \DP_OP_379J1_125_371/n196 ), .CI(\DP_OP_379J1_125_371/n43 ), .CO(
        \DP_OP_379J1_125_371/n42 ), .S(N109) );
  FA1D0BWP \DP_OP_379J1_125_371/U54  ( .A(\DP_OP_379J1_125_371/n131 ), .B(
        \DP_OP_379J1_125_371/n135 ), .CI(\DP_OP_379J1_125_371/n42 ), .CO(
        \DP_OP_379J1_125_371/n41 ), .S(N110) );
  FA1D0BWP \DP_OP_379J1_125_371/U53  ( .A(\DP_OP_379J1_125_371/n129 ), .B(
        \DP_OP_379J1_125_371/n130 ), .CI(\DP_OP_379J1_125_371/n41 ), .CO(
        \DP_OP_379J1_125_371/n40 ), .S(N111) );
  FA1D0BWP \DP_OP_379J1_125_371/U52  ( .A(\DP_OP_379J1_125_371/n125 ), .B(
        \DP_OP_379J1_125_371/n128 ), .CI(\DP_OP_379J1_125_371/n40 ), .CO(
        \DP_OP_379J1_125_371/n39 ), .S(N112) );
  FA1D0BWP \DP_OP_379J1_125_371/U51  ( .A(\DP_OP_379J1_125_371/n123 ), .B(
        \DP_OP_379J1_125_371/n124 ), .CI(\DP_OP_379J1_125_371/n39 ), .CO(
        \DP_OP_379J1_125_371/n38 ), .S(N113) );
  FA1D0BWP \DP_OP_379J1_125_371/U50  ( .A(\DP_OP_379J1_125_371/n122 ), .B(
        \DP_OP_379J1_125_371/n118 ), .CI(\DP_OP_379J1_125_371/n38 ), .CO(
        \DP_OP_379J1_125_371/n37 ), .S(N114) );
  FA1D0BWP \DP_OP_379J1_125_371/U49  ( .A(\DP_OP_379J1_125_371/n113 ), .B(
        \DP_OP_379J1_125_371/n117 ), .CI(\DP_OP_379J1_125_371/n37 ), .CO(
        \DP_OP_379J1_125_371/n36 ), .S(N115) );
  FA1D0BWP \DP_OP_379J1_125_371/U48  ( .A(\DP_OP_379J1_125_371/n106 ), .B(
        \DP_OP_379J1_125_371/n112 ), .CI(\DP_OP_379J1_125_371/n36 ), .CO(
        \DP_OP_379J1_125_371/n35 ), .S(N116) );
  FA1D0BWP \DP_OP_379J1_125_371/U47  ( .A(\DP_OP_379J1_125_371/n100 ), .B(
        \DP_OP_379J1_125_371/n105 ), .CI(\DP_OP_379J1_125_371/n35 ), .CO(
        \DP_OP_379J1_125_371/n34 ), .S(N117) );
  FA1D0BWP \DP_OP_379J1_125_371/U46  ( .A(\DP_OP_379J1_125_371/n94 ), .B(
        \DP_OP_379J1_125_371/n99 ), .CI(\DP_OP_379J1_125_371/n34 ), .CO(
        \DP_OP_379J1_125_371/n33 ), .S(N118) );
  FA1D0BWP \DP_OP_379J1_125_371/U45  ( .A(\DP_OP_379J1_125_371/n87 ), .B(
        \DP_OP_379J1_125_371/n93 ), .CI(\DP_OP_379J1_125_371/n33 ), .CO(
        \DP_OP_379J1_125_371/n32 ), .S(N119) );
  FA1D0BWP \DP_OP_379J1_125_371/U44  ( .A(\DP_OP_379J1_125_371/n79 ), .B(
        \DP_OP_379J1_125_371/n86 ), .CI(\DP_OP_379J1_125_371/n32 ), .CO(
        \DP_OP_379J1_125_371/n31 ), .S(N120) );
  FA1D0BWP \DP_OP_379J1_125_371/U43  ( .A(\DP_OP_379J1_125_371/n78 ), .B(
        \DP_OP_379J1_125_371/n73 ), .CI(\DP_OP_379J1_125_371/n31 ), .CO(
        \DP_OP_379J1_125_371/n30 ), .S(N121) );
  FA1D0BWP \DP_OP_379J1_125_371/U42  ( .A(\DP_OP_379J1_125_371/n72 ), .B(
        \DP_OP_379J1_125_371/n66 ), .CI(\DP_OP_379J1_125_371/n30 ), .CO(
        \DP_OP_379J1_125_371/n29 ), .S(N122) );
  FA1D0BWP \DP_OP_379J1_125_371/U41  ( .A(\DP_OP_379J1_125_371/n65 ), .B(
        \DP_OP_379J1_125_371/n61 ), .CI(\DP_OP_379J1_125_371/n29 ), .CO(
        \DP_OP_379J1_125_371/n28 ), .S(N123) );
  FA1D0BWP \DP_OP_379J1_125_371/U40  ( .A(\DP_OP_379J1_125_371/n60 ), .B(
        \DP_OP_379J1_125_371/n56 ), .CI(\DP_OP_379J1_125_371/n28 ), .CO(
        \DP_OP_379J1_125_371/n27 ), .S(N124) );
  FA1D0BWP \DP_OP_379J1_125_371/U39  ( .A(\DP_OP_379J1_125_371/n55 ), .B(
        \DP_OP_379J1_125_371/n53 ), .CI(\DP_OP_379J1_125_371/n27 ), .CO(
        \DP_OP_379J1_125_371/n26 ), .S(N125) );
  FA1D0BWP \DP_OP_379J1_125_371/U38  ( .A(\DP_OP_379J1_125_371/n52 ), .B(
        \DP_OP_379J1_125_371/n48 ), .CI(\DP_OP_379J1_125_371/n26 ), .CO(
        \DP_OP_379J1_125_371/n25 ), .S(N126) );
  AO22D1BWP \DP_OP_379J1_125_371/U32  ( .A1(N117), .A2(
        \DP_OP_379J1_125_371/I5 ), .B1(\DP_OP_379J1_125_371/I4 ), .B2(N1782), 
        .Z(\DP_OP_379J1_125_371/n9 ) );
  AO22D1BWP \DP_OP_379J1_125_371/U31  ( .A1(N118), .A2(
        \DP_OP_379J1_125_371/I5 ), .B1(\DP_OP_379J1_125_371/I4 ), .B2(N1783), 
        .Z(\DP_OP_379J1_125_371/n335 ) );
  AO22D1BWP \DP_OP_379J1_125_371/U30  ( .A1(N119), .A2(
        \DP_OP_379J1_125_371/I5 ), .B1(\DP_OP_379J1_125_371/I4 ), .B2(N1784), 
        .Z(\DP_OP_379J1_125_371/n336 ) );
  AO22D1BWP \DP_OP_379J1_125_371/U29  ( .A1(N120), .A2(
        \DP_OP_379J1_125_371/I5 ), .B1(\DP_OP_379J1_125_371/I4 ), .B2(N1785), 
        .Z(\DP_OP_379J1_125_371/n337 ) );
  AO22D1BWP \DP_OP_379J1_125_371/U28  ( .A1(N121), .A2(
        \DP_OP_379J1_125_371/I5 ), .B1(\DP_OP_379J1_125_371/I4 ), .B2(N1786), 
        .Z(\DP_OP_379J1_125_371/n338 ) );
  AO22D1BWP \DP_OP_379J1_125_371/U27  ( .A1(N122), .A2(
        \DP_OP_379J1_125_371/I5 ), .B1(\DP_OP_379J1_125_371/I4 ), .B2(N1787), 
        .Z(\DP_OP_379J1_125_371/n339 ) );
  AO22D1BWP \DP_OP_379J1_125_371/U26  ( .A1(N123), .A2(
        \DP_OP_379J1_125_371/I5 ), .B1(\DP_OP_379J1_125_371/I4 ), .B2(N1788), 
        .Z(\DP_OP_379J1_125_371/n340 ) );
  AO22D1BWP \DP_OP_379J1_125_371/U25  ( .A1(N124), .A2(
        \DP_OP_379J1_125_371/I5 ), .B1(\DP_OP_379J1_125_371/I4 ), .B2(N1789), 
        .Z(\DP_OP_379J1_125_371/n341 ) );
  AO22D1BWP \DP_OP_379J1_125_371/U24  ( .A1(N125), .A2(
        \DP_OP_379J1_125_371/I5 ), .B1(\DP_OP_379J1_125_371/I4 ), .B2(N1790), 
        .Z(\DP_OP_379J1_125_371/n342 ) );
  OAI22D1BWP \DP_OP_379J1_125_371/U95  ( .A1(\DP_OP_379J1_125_371/n319 ), .A2(
        n533), .B1(\DP_OP_379J1_125_371/n325 ), .B2(n534), .ZN(
        \DP_OP_379J1_125_371/n49 ) );
  FA1D0BWP \DP_OP_379J1_125_371/U58  ( .A(\DP_OP_379J1_125_371/n138 ), .B(
        \DP_OP_379J1_125_371/n49 ), .CI(\DP_OP_379J1_125_371/n145 ), .CO(
        \DP_OP_379J1_125_371/n45 ), .S(\DP_OP_379J1_125_371/n46 ) );
  INR2D1BWP \DP_OP_379J1_125_371/U233  ( .A1(B[0]), .B1(n536), .ZN(N107) );
  FA1D0BWP \DP_OP_379J1_125_371/U37  ( .A(\DP_OP_379J1_125_371/n47 ), .B(
        \DP_OP_379J1_125_371/n46 ), .CI(\DP_OP_379J1_125_371/n25 ), .CO(
        \DP_OP_379J1_125_371/n24 ), .S(N127) );
  CKND2D0BWP \DP_OP_379J1_125_371/U278  ( .A1(\DP_OP_379J1_125_371/n325 ), 
        .A2(N92), .ZN(\DP_OP_379J1_125_371/n319 ) );
  HA1D0BWP \DP_OP_379J1_125_371/U90  ( .A(\DP_OP_379J1_125_371/n134 ), .B(
        \DP_OP_379J1_125_371/n182 ), .CO(\DP_OP_379J1_125_371/n126 ), .S(
        \DP_OP_379J1_125_371/n127 ) );
  HA1D0BWP \DP_OP_379J1_125_371/U92  ( .A(\DP_OP_379J1_125_371/n195 ), .B(
        \DP_OP_379J1_125_371/n206 ), .CO(\DP_OP_379J1_125_371/n130 ), .S(
        \DP_OP_379J1_125_371/n131 ) );
  HA1D0BWP \DP_OP_379J1_125_371/U56  ( .A(\DP_OP_379J1_125_371/n208 ), .B(
        \DP_OP_379J1_125_371/n136 ), .CO(\DP_OP_379J1_125_371/n43 ), .S(N108)
         );
  HA1D0BWP \DP_OP_379J1_125_371/U21  ( .A(N119), .B(N118), .CO(
        \DP_OP_379J1_125_371/n19 ), .S(N141) );
  HA1D0BWP \DP_OP_379J1_125_371/U20  ( .A(N120), .B(\DP_OP_379J1_125_371/n19 ), 
        .CO(\DP_OP_379J1_125_371/n18 ), .S(N142) );
  HA1D0BWP \DP_OP_379J1_125_371/U19  ( .A(N121), .B(\DP_OP_379J1_125_371/n18 ), 
        .CO(\DP_OP_379J1_125_371/n17 ), .S(N143) );
  HA1D0BWP \DP_OP_379J1_125_371/U18  ( .A(N122), .B(\DP_OP_379J1_125_371/n17 ), 
        .CO(\DP_OP_379J1_125_371/n16 ), .S(N144) );
  HA1D0BWP \DP_OP_379J1_125_371/U17  ( .A(N123), .B(\DP_OP_379J1_125_371/n16 ), 
        .CO(\DP_OP_379J1_125_371/n15 ), .S(N145) );
  HA1D0BWP \DP_OP_379J1_125_371/U16  ( .A(N124), .B(\DP_OP_379J1_125_371/n15 ), 
        .CO(\DP_OP_379J1_125_371/n14 ), .S(N146) );
  HA1D0BWP \DP_OP_379J1_125_371/U15  ( .A(N125), .B(\DP_OP_379J1_125_371/n14 ), 
        .CO(\DP_OP_379J1_125_371/n13 ), .S(N147) );
  HA1D0BWP \DP_OP_379J1_125_371/U14  ( .A(N126), .B(\DP_OP_379J1_125_371/n13 ), 
        .CO(\DP_OP_379J1_125_371/n12 ), .S(N148) );
  HA1D0BWP \DP_OP_379J1_125_371/U13  ( .A(N127), .B(\DP_OP_379J1_125_371/n12 ), 
        .CO(\DP_OP_379J1_125_371/n11 ), .S(N149) );
  HA1D0BWP \DP_OP_379J1_125_371/U12  ( .A(N1940), .B(\DP_OP_379J1_125_371/n11 ), .CO(\DP_OP_379J1_125_371/n10 ), .S(N150) );
  HA1D0BWP \DP_OP_379J1_125_371/U9  ( .A(\DP_OP_379J1_125_371/n335 ), .B(
        \DP_OP_379J1_125_371/n9 ), .CO(\DP_OP_379J1_125_371/n8 ), .S(
        \C148/DATA4_1 ) );
  HA1D0BWP \DP_OP_379J1_125_371/U8  ( .A(\DP_OP_379J1_125_371/n336 ), .B(
        \DP_OP_379J1_125_371/n8 ), .CO(\DP_OP_379J1_125_371/n7 ), .S(
        \C148/DATA4_2 ) );
  HA1D0BWP \DP_OP_379J1_125_371/U7  ( .A(\DP_OP_379J1_125_371/n337 ), .B(
        \DP_OP_379J1_125_371/n7 ), .CO(\DP_OP_379J1_125_371/n6 ), .S(
        \C148/DATA4_3 ) );
  HA1D0BWP \DP_OP_379J1_125_371/U6  ( .A(\DP_OP_379J1_125_371/n338 ), .B(
        \DP_OP_379J1_125_371/n6 ), .CO(\DP_OP_379J1_125_371/n5 ), .S(
        \C148/DATA4_4 ) );
  HA1D0BWP \DP_OP_379J1_125_371/U5  ( .A(\DP_OP_379J1_125_371/n339 ), .B(
        \DP_OP_379J1_125_371/n5 ), .CO(\DP_OP_379J1_125_371/n4 ), .S(
        \C148/DATA4_5 ) );
  HA1D0BWP \DP_OP_379J1_125_371/U4  ( .A(\DP_OP_379J1_125_371/n340 ), .B(
        \DP_OP_379J1_125_371/n4 ), .CO(\DP_OP_379J1_125_371/n3 ), .S(
        \C148/DATA4_6 ) );
  HA1D0BWP \DP_OP_379J1_125_371/U3  ( .A(\DP_OP_379J1_125_371/n341 ), .B(
        \DP_OP_379J1_125_371/n3 ), .CO(\DP_OP_379J1_125_371/n2 ), .S(
        \C148/DATA4_7 ) );
  HA1D0BWP \DP_OP_379J1_125_371/U2  ( .A(\DP_OP_379J1_125_371/n342 ), .B(
        \DP_OP_379J1_125_371/n2 ), .CO(\DP_OP_379J1_125_371/n1 ), .S(
        \C148/DATA4_8 ) );
  CKND0BWP \DP_OP_379J1_125_371/U10  ( .I(\DP_OP_379J1_125_371/n9 ), .ZN(
        \C148/DATA4_0 ) );
  HA1D0BWP \DP_OP_379J1_125_371/U83  ( .A(\DP_OP_379J1_125_371/n132 ), .B(
        \DP_OP_379J1_125_371/n156 ), .CO(\DP_OP_379J1_125_371/n109 ), .S(
        \DP_OP_379J1_125_371/n110 ) );
  HA1D0BWP \DP_OP_379J1_125_371/U87  ( .A(\DP_OP_379J1_125_371/n133 ), .B(
        \DP_OP_379J1_125_371/n169 ), .CO(\DP_OP_379J1_125_371/n119 ), .S(
        \DP_OP_379J1_125_371/n120 ) );
  INVD1BWP U519 ( .I(n941), .ZN(n766) );
  XNR2D1BWP U520 ( .A1(A[2]), .A2(A[1]), .ZN(\DP_OP_379J1_125_371/n329 ) );
  XNR2D1BWP U521 ( .A1(A[4]), .A2(A[3]), .ZN(\DP_OP_379J1_125_371/n328 ) );
  XNR2D1BWP U522 ( .A1(A[6]), .A2(A[5]), .ZN(\DP_OP_379J1_125_371/n327 ) );
  INVD1BWP U523 ( .I(A[0]), .ZN(n536) );
  OAI31D1BWP U524 ( .A1(n1337), .A2(n1338), .A3(n1239), .B(n1238), .ZN(n1325)
         );
  INVD1BWP U525 ( .I(B[10]), .ZN(n765) );
  XNR2D1BWP U526 ( .A1(A[8]), .A2(A[7]), .ZN(\DP_OP_379J1_125_371/n326 ) );
  XNR2D1BWP U527 ( .A1(N92), .A2(A[9]), .ZN(\DP_OP_379J1_125_371/n325 ) );
  NR2XD1BWP U528 ( .A1(n746), .A2(n1325), .ZN(n751) );
  OAI222D0BWP U529 ( .A1(n1115), .A2(n1118), .B1(n758), .B2(n1117), .C1(n1116), 
        .C2(n1112), .ZN(n1175) );
  CKND0BWP U530 ( .I(n1252), .ZN(n446) );
  NR2D0BWP U531 ( .A1(n1253), .A2(n1256), .ZN(n447) );
  MUX2ND0BWP U532 ( .I0(n1252), .I1(n446), .S(n447), .ZN(n1273) );
  IAO21D0BWP U533 ( .A1(n1227), .A2(n1231), .B(n1222), .ZN(n1220) );
  CKND0BWP U534 ( .I(n782), .ZN(n448) );
  AO21D0BWP U535 ( .A1(N125), .A2(n448), .B(n549), .Z(n550) );
  OAI31D0BWP U536 ( .A1(n698), .A2(n855), .A3(n854), .B(n607), .ZN(n898) );
  MOAI22D0BWP U537 ( .A1(n735), .A2(n666), .B1(\C148/DATA4_4 ), .B2(n719), 
        .ZN(n449) );
  OAI22D0BWP U538 ( .A1(n736), .A2(n668), .B1(n667), .B2(n673), .ZN(n450) );
  AO211D0BWP U539 ( .A1(n712), .A2(N1786), .B(n449), .C(n450), .Z(N1850) );
  CKND0BWP U540 ( .I(n1104), .ZN(n451) );
  INR2D0BWP U541 ( .A1(n1103), .B1(n1119), .ZN(n452) );
  MUX2ND0BWP U542 ( .I0(n1104), .I1(n451), .S(n452), .ZN(n1135) );
  IND2D0BWP U543 ( .A1(n785), .B1(n783), .ZN(n790) );
  CKND0BWP U544 ( .I(n925), .ZN(n453) );
  MUX2ND0BWP U545 ( .I0(n453), .I1(n925), .S(n926), .ZN(n454) );
  CKND0BWP U546 ( .I(n927), .ZN(n455) );
  AOI211D0BWP U547 ( .A1(n934), .A2(n956), .B(n928), .C(n931), .ZN(n456) );
  OAI211D0BWP U548 ( .A1(n923), .A2(n919), .B(n930), .C(n456), .ZN(n457) );
  OAI31D0BWP U549 ( .A1(n454), .A2(n455), .A3(n457), .B(n911), .ZN(n939) );
  CKND2D0BWP U550 ( .A1(A[2]), .A2(A[3]), .ZN(n458) );
  OAI211D0BWP U551 ( .A1(A[2]), .A2(A[3]), .B(\DP_OP_379J1_125_371/n329 ), .C(
        n458), .ZN(\DP_OP_379J1_125_371/n323 ) );
  CKND0BWP U552 ( .I(n1216), .ZN(n459) );
  OAI22D0BWP U553 ( .A1(n459), .A2(n1215), .B1(n1231), .B2(n1227), .ZN(n460)
         );
  AOI221D0BWP U554 ( .A1(n459), .A2(n1215), .B1(n1227), .B2(n1231), .C(n460), 
        .ZN(n461) );
  ND3D0BWP U555 ( .A1(n1223), .A2(n1226), .A3(n1207), .ZN(n462) );
  AOI211D0BWP U556 ( .A1(n1205), .A2(n1206), .B(n1220), .C(n462), .ZN(n463) );
  AOI211D0BWP U557 ( .A1(n461), .A2(n463), .B(n1208), .C(n1209), .ZN(n1232) );
  IND2D0BWP U558 ( .A1(n550), .B1(n551), .ZN(n913) );
  MOAI22D0BWP U559 ( .A1(n735), .A2(n668), .B1(\C148/DATA4_5 ), .B2(n719), 
        .ZN(n464) );
  OAI22D0BWP U560 ( .A1(n736), .A2(n670), .B1(n669), .B2(n673), .ZN(n465) );
  AO211D0BWP U561 ( .A1(n712), .A2(N1787), .B(n464), .C(n465), .Z(N1851) );
  CKND0BWP U562 ( .I(n1135), .ZN(n466) );
  NR2D0BWP U563 ( .A1(n1137), .A2(n1136), .ZN(n467) );
  MUX2ND0BWP U564 ( .I0(n1135), .I1(n466), .S(n467), .ZN(n1161) );
  AOI22D0BWP U565 ( .A1(n1084), .A2(n1083), .B1(n1081), .B2(n1082), .ZN(n468)
         );
  OA21D0BWP U566 ( .A1(n1050), .A2(n1049), .B(n468), .Z(n1115) );
  ND4D0BWP U567 ( .A1(n592), .A2(n599), .A3(n596), .A4(n600), .ZN(n469) );
  NR3D0BWP U568 ( .A1(n607), .A2(n603), .A3(n469), .ZN(n470) );
  AOI21D0BWP U569 ( .A1(n753), .A2(n470), .B(n782), .ZN(n551) );
  NR2D0BWP U570 ( .A1(n1025), .A2(n1028), .ZN(n471) );
  CKND2D0BWP U571 ( .A1(n997), .A2(n996), .ZN(n472) );
  OAI211D0BWP U572 ( .A1(n997), .A2(n996), .B(n1034), .C(n472), .ZN(n473) );
  NR4D0BWP U573 ( .A1(n1016), .A2(n1019), .A3(n471), .A4(n473), .ZN(n474) );
  AOI31D0BWP U574 ( .A1(n1032), .A2(n1027), .A3(n474), .B(n1005), .ZN(n1040)
         );
  CKND2D0BWP U575 ( .A1(A[4]), .A2(A[5]), .ZN(n475) );
  OAI211D0BWP U576 ( .A1(A[4]), .A2(A[5]), .B(\DP_OP_379J1_125_371/n328 ), .C(
        n475), .ZN(\DP_OP_379J1_125_371/n322 ) );
  INR2D0BWP U577 ( .A1(n1258), .B1(n1269), .ZN(n476) );
  NR4D0BWP U578 ( .A1(n1246), .A2(n1251), .A3(n1260), .A4(n476), .ZN(n477) );
  OAI211D0BWP U579 ( .A1(n1252), .A2(n1217), .B(n477), .C(n1254), .ZN(n478) );
  AOI21D0BWP U580 ( .A1(n1252), .A2(n1217), .B(n478), .ZN(n479) );
  MAOI22D0BWP U581 ( .A1(n1244), .A2(n1242), .B1(n1244), .B2(n1242), .ZN(n480)
         );
  IOA21D0BWP U582 ( .A1(n480), .A2(n479), .B(n1232), .ZN(n1240) );
  MOAI22D0BWP U583 ( .A1(n735), .A2(n670), .B1(\C148/DATA4_6 ), .B2(n719), 
        .ZN(n481) );
  OAI22D0BWP U584 ( .A1(n736), .A2(n672), .B1(n673), .B2(n671), .ZN(n482) );
  AO211D0BWP U585 ( .A1(n712), .A2(N1788), .B(n481), .C(n482), .Z(N1852) );
  CKND0BWP U586 ( .I(n899), .ZN(n483) );
  NR2D0BWP U587 ( .A1(n1315), .A2(n900), .ZN(n484) );
  MUX2ND0BWP U588 ( .I0(n899), .I1(n483), .S(n484), .ZN(n931) );
  NR2D0BWP U589 ( .A1(n1091), .A2(n1095), .ZN(n485) );
  OAI211D0BWP U590 ( .A1(n1101), .A2(n1103), .B(n1104), .C(n485), .ZN(n486) );
  AOI211D0BWP U591 ( .A1(n1069), .A2(n1070), .B(n1105), .C(n486), .ZN(n487) );
  OAI21D0BWP U592 ( .A1(n1069), .A2(n1070), .B(n487), .ZN(n488) );
  IAO21D0BWP U593 ( .A1(n1094), .A2(n488), .B(n1076), .ZN(n1111) );
  CKND0BWP U594 ( .I(n1198), .ZN(n489) );
  NR2D0BWP U595 ( .A1(n1200), .A2(n1199), .ZN(n490) );
  MUX2ND0BWP U596 ( .I0(n1198), .I1(n489), .S(n490), .ZN(n1227) );
  NR3D0BWP U597 ( .A1(n1270), .A2(n1282), .A3(n1273), .ZN(n491) );
  CKND0BWP U598 ( .I(n1291), .ZN(n492) );
  OAI22D0BWP U599 ( .A1(n492), .A2(n1261), .B1(n1266), .B2(n1267), .ZN(n493)
         );
  AOI221D0BWP U600 ( .A1(n492), .A2(n1261), .B1(n1267), .B2(n1266), .C(n493), 
        .ZN(n494) );
  ND4D0BWP U601 ( .A1(n1264), .A2(n1268), .A3(n491), .A4(n494), .ZN(n495) );
  ND3D0BWP U602 ( .A1(n1320), .A2(n1262), .A3(n495), .ZN(n1305) );
  INR3D0BWP U603 ( .A1(n795), .B1(n800), .B2(n794), .ZN(n496) );
  IND4D0BWP U604 ( .A1(n789), .B1(n803), .B2(n496), .B3(n798), .ZN(n497) );
  OAI31D0BWP U605 ( .A1(n607), .A2(n790), .A3(n497), .B(n551), .ZN(n806) );
  CKND2D0BWP U606 ( .A1(A[8]), .A2(A[9]), .ZN(n498) );
  OAI211D0BWP U607 ( .A1(A[8]), .A2(A[9]), .B(\DP_OP_379J1_125_371/n326 ), .C(
        n498), .ZN(\DP_OP_379J1_125_371/n320 ) );
  INR2D0BWP U608 ( .A1(n587), .B1(n1053), .ZN(N1783) );
  MOAI22D0BWP U609 ( .A1(n735), .A2(n672), .B1(\C148/DATA4_7 ), .B2(n719), 
        .ZN(n499) );
  OAI22D0BWP U610 ( .A1(n736), .A2(n678), .B1(n673), .B2(n674), .ZN(n500) );
  AO211D0BWP U611 ( .A1(n712), .A2(N1789), .B(n499), .C(n500), .Z(N1853) );
  IOA21D0BWP U612 ( .A1(n1260), .A2(n1259), .B(n1270), .ZN(n1271) );
  CKND0BWP U613 ( .I(n1315), .ZN(n501) );
  AOI31D0BWP U614 ( .A1(n899), .A2(n897), .A3(n501), .B(n898), .ZN(n956) );
  CKND0BWP U615 ( .I(n824), .ZN(n502) );
  IND3D0BWP U616 ( .A1(n1313), .B1(n826), .B2(n825), .ZN(n503) );
  MUX2ND0BWP U617 ( .I0(n502), .I1(n824), .S(n503), .ZN(n834) );
  CKND0BWP U618 ( .I(n857), .ZN(n504) );
  OAI32D0BWP U619 ( .A1(n504), .A2(n698), .A3(n856), .B1(n858), .B2(n504), 
        .ZN(n879) );
  CKND0BWP U620 ( .I(n1129), .ZN(n505) );
  MUX2ND0BWP U621 ( .I0(n505), .I1(n1129), .S(n1128), .ZN(n506) );
  CKND0BWP U622 ( .I(n1110), .ZN(n507) );
  AOI211D0BWP U623 ( .A1(n1137), .A2(n1159), .B(n1131), .C(n1135), .ZN(n508)
         );
  OAI211D0BWP U624 ( .A1(n1122), .A2(n1126), .B(n1134), .C(n508), .ZN(n509) );
  OAI31D0BWP U625 ( .A1(n506), .A2(n507), .A3(n509), .B(n1111), .ZN(n1141) );
  AO21D0BWP U626 ( .A1(n1294), .A2(n1291), .B(n1269), .Z(n1268) );
  CKND2D0BWP U627 ( .A1(A[0]), .A2(A[1]), .ZN(n510) );
  OAI211D0BWP U628 ( .A1(A[0]), .A2(A[1]), .B(n536), .C(n510), .ZN(
        \DP_OP_379J1_125_371/n324 ) );
  NR4D0BWP U629 ( .A1(A[14]), .A2(A[10]), .A3(A[11]), .A4(A[13]), .ZN(n511) );
  IND2D0BWP U630 ( .A1(A[12]), .B1(n511), .ZN(N92) );
  NR4D0BWP U631 ( .A1(B[12]), .A2(B[11]), .A3(B[13]), .A4(B[10]), .ZN(n512) );
  CKND2D0BWP U632 ( .A1(n764), .A2(n512), .ZN(N93) );
  CKND0BWP U633 ( .I(n1116), .ZN(n513) );
  OA221D0BWP U634 ( .A1(n1116), .A2(n587), .B1(n513), .B2(n586), .C(n1173), 
        .Z(N1784) );
  AOI22D0BWP U635 ( .A1(N126), .A2(n711), .B1(n730), .B2(N150), .ZN(n514) );
  AO22D0BWP U636 ( .A1(\DP_OP_379J1_125_371/I4 ), .A2(N1791), .B1(
        \DP_OP_379J1_125_371/I5 ), .B2(N126), .Z(n515) );
  CKND2D0BWP U637 ( .A1(\DP_OP_379J1_125_371/n1 ), .A2(n515), .ZN(n516) );
  OAI211D0BWP U638 ( .A1(\DP_OP_379J1_125_371/n1 ), .A2(n515), .B(n719), .C(
        n516), .ZN(n517) );
  OAI211D0BWP U639 ( .A1(n735), .A2(n680), .B(n514), .C(n517), .ZN(n518) );
  AO21D0BWP U640 ( .A1(n712), .A2(N1791), .B(n518), .Z(N1855) );
  NR2D0BWP U641 ( .A1(n889), .A2(n901), .ZN(n519) );
  OAI211D0BWP U642 ( .A1(n898), .A2(n897), .B(n899), .C(n519), .ZN(n520) );
  AOI211D0BWP U643 ( .A1(n890), .A2(n893), .B(n904), .C(n520), .ZN(n521) );
  OAI21D0BWP U644 ( .A1(n890), .A2(n893), .B(n521), .ZN(n522) );
  IAO21D0BWP U645 ( .A1(n896), .A2(n522), .B(n909), .ZN(n911) );
  CKND2D0BWP U646 ( .A1(A[6]), .A2(A[7]), .ZN(n523) );
  OAI211D0BWP U647 ( .A1(A[6]), .A2(A[7]), .B(\DP_OP_379J1_125_371/n327 ), .C(
        n523), .ZN(\DP_OP_379J1_125_371/n321 ) );
  IAO21D0BWP U648 ( .A1(n1337), .A2(n1328), .B(n774), .ZN(n1329) );
  IND2D0BWP U649 ( .A1(n806), .B1(n552), .ZN(n1313) );
  INR2D0BWP U650 ( .A1(n585), .B1(n1176), .ZN(N1785) );
  INR2D0BWP U651 ( .A1(n579), .B1(n1221), .ZN(N1789) );
  INR2D0BWP U652 ( .A1(n638), .B1(n756), .ZN(N1791) );
  INR2D0BWP U653 ( .A1(N107), .B1(n751), .ZN(N1919) );
  NR2D0BWP U654 ( .A1(\DP_OP_379J1_125_371/n319 ), .A2(n535), .ZN(n524) );
  XNR3D0BWP U655 ( .A1(\DP_OP_379J1_125_371/n45 ), .A2(n524), .A3(
        \DP_OP_379J1_125_371/n24 ), .ZN(N1940) );
  ND2D1BWP U656 ( .A1(n1346), .A2(n1349), .ZN(N78) );
  INVD1BWP U657 ( .I(n1313), .ZN(n761) );
  CKND2D0BWP U658 ( .A1(N115), .A2(n546), .ZN(n705) );
  CKND2D0BWP U659 ( .A1(N107), .A2(n683), .ZN(n681) );
  CKND0BWP U660 ( .I(N1791), .ZN(n707) );
  CKND0BWP U661 ( .I(n1310), .ZN(n1311) );
  CKND2D0BWP U662 ( .A1(n751), .A2(n941), .ZN(n701) );
  CKND2D0BWP U663 ( .A1(N112), .A2(n546), .ZN(n695) );
  CKND0BWP U664 ( .I(n697), .ZN(n696) );
  CKND0BWP U665 ( .I(n751), .ZN(n546) );
  CKND0BWP U666 ( .I(\DP_OP_379J1_125_371/n83 ), .ZN(n542) );
  CKND0BWP U667 ( .I(\DP_OP_379J1_125_371/n57 ), .ZN(n544) );
  CKND0BWP U668 ( .I(\DP_OP_379J1_125_371/n69 ), .ZN(n543) );
  CKND0BWP U669 ( .I(B[4]), .ZN(n529) );
  CKND0BWP U670 ( .I(B[3]), .ZN(n528) );
  CKND0BWP U671 ( .I(B[0]), .ZN(n525) );
  CKND0BWP U672 ( .I(B[5]), .ZN(n530) );
  CKND0BWP U673 ( .I(B[2]), .ZN(n527) );
  CKND0BWP U674 ( .I(B[1]), .ZN(n526) );
  CKND0BWP U675 ( .I(A[7]), .ZN(n540) );
  CKND0BWP U676 ( .I(B[6]), .ZN(n531) );
  CKND0BWP U677 ( .I(B[7]), .ZN(n532) );
  CKND2D0BWP U678 ( .A1(A[15]), .A2(n1346), .ZN(n1348) );
  CKND0BWP U679 ( .I(A[15]), .ZN(n1350) );
  CKND2D0BWP U680 ( .A1(n712), .A2(N1782), .ZN(n716) );
  MAOI22D0BWP U681 ( .A1(N117), .A2(n711), .B1(n710), .B2(n736), .ZN(n717) );
  CKND0BWP U682 ( .I(n711), .ZN(n673) );
  CKND2D0BWP U683 ( .A1(n1326), .A2(n741), .ZN(n723) );
  CKND0BWP U684 ( .I(n1291), .ZN(n1293) );
  CKND2D0BWP U685 ( .A1(n745), .A2(n727), .ZN(prod[11]) );
  CKND0BWP U686 ( .I(n1287), .ZN(n1303) );
  CKAN2D0BWP U687 ( .A1(n1332), .A2(n1331), .Z(n1336) );
  OR2XD1BWP U688 ( .A1(n1301), .A2(n1300), .Z(n1331) );
  CKND2D0BWP U689 ( .A1(n1337), .A2(n731), .ZN(n728) );
  CKND0BWP U690 ( .I(n742), .ZN(n729) );
  CKND0BWP U691 ( .I(n1338), .ZN(n1340) );
  CKND0BWP U692 ( .I(n1307), .ZN(n1342) );
  CKND2D0BWP U693 ( .A1(n1301), .A2(n1300), .ZN(n1332) );
  CKND2D0BWP U694 ( .A1(n1278), .A2(n1285), .ZN(n1287) );
  CKND0BWP U695 ( .I(n1286), .ZN(n1280) );
  CKND2D0BWP U696 ( .A1(n1286), .A2(n1285), .ZN(n1288) );
  CKND0BWP U697 ( .I(n1281), .ZN(n1285) );
  CKND2D0BWP U698 ( .A1(n756), .A2(n1270), .ZN(n1272) );
  CKND2D0BWP U699 ( .A1(n756), .A2(n1263), .ZN(n1274) );
  CKND0BWP U700 ( .I(n1273), .ZN(n1276) );
  CKND0BWP U701 ( .I(n1261), .ZN(n1294) );
  CKND0BWP U702 ( .I(n1254), .ZN(n1257) );
  CKND0BWP U703 ( .I(n1240), .ZN(n1262) );
  CKND2D0BWP U704 ( .A1(n735), .A2(n736), .ZN(n742) );
  CKND0BWP U705 ( .I(n741), .ZN(n743) );
  CKND0BWP U706 ( .I(n720), .ZN(n721) );
  CKND2D0BWP U707 ( .A1(n714), .A2(N1940), .ZN(n720) );
  CKND0BWP U708 ( .I(n750), .ZN(n722) );
  CKND0BWP U709 ( .I(n1299), .ZN(n1345) );
  CKND0BWP U710 ( .I(n756), .ZN(n1295) );
  CKND0BWP U711 ( .I(n1227), .ZN(n1230) );
  CKND2D0BWP U712 ( .A1(n1242), .A2(n1244), .ZN(n1258) );
  CKND0BWP U713 ( .I(n1232), .ZN(n1235) );
  CKND0BWP U714 ( .I(n1242), .ZN(n1245) );
  CKND2D0BWP U715 ( .A1(n1264), .A2(n1263), .ZN(n1266) );
  CKND2D0BWP U716 ( .A1(n1251), .A2(n1250), .ZN(n1259) );
  CKND0BWP U717 ( .I(n1250), .ZN(n1256) );
  CKND0BWP U718 ( .I(n1246), .ZN(n1248) );
  CKND2D0BWP U719 ( .A1(n1252), .A2(n1217), .ZN(n1249) );
  CKND0BWP U720 ( .I(n1253), .ZN(n1217) );
  CKND2D0BWP U721 ( .A1(n1251), .A2(n1226), .ZN(n1253) );
  CKND0BWP U722 ( .I(n1221), .ZN(n1229) );
  CKND2D0BWP U723 ( .A1(n1211), .A2(n1221), .ZN(n1224) );
  CKND0BWP U724 ( .I(n736), .ZN(n730) );
  CKND2D0BWP U725 ( .A1(\C148/DATA4_8 ), .A2(n719), .ZN(n676) );
  MAOI22D0BWP U726 ( .A1(N125), .A2(n711), .B1(n680), .B2(n736), .ZN(n677) );
  CKND2D0BWP U727 ( .A1(N1940), .A2(n648), .ZN(n736) );
  CKND0BWP U728 ( .I(n649), .ZN(n650) );
  CKND2D0BWP U729 ( .A1(N116), .A2(N117), .ZN(n649) );
  CKND2D0BWP U730 ( .A1(N127), .A2(n646), .ZN(n741) );
  CKND0BWP U731 ( .I(n731), .ZN(n735) );
  CKND0BWP U732 ( .I(\DP_OP_379J1_125_371/n10 ), .ZN(n645) );
  CKND0BWP U733 ( .I(n647), .ZN(n675) );
  CKND2D0BWP U734 ( .A1(N117), .A2(N118), .ZN(n647) );
  CKAN2D0BWP U735 ( .A1(n1232), .A2(n1233), .Z(n1250) );
  CKND0BWP U736 ( .I(n1210), .ZN(n1188) );
  CKND2D0BWP U737 ( .A1(n1201), .A2(n755), .ZN(n1204) );
  XNR2D1BWP U738 ( .A1(n1194), .A2(n1205), .ZN(n1219) );
  CKND2D0BWP U739 ( .A1(n1207), .A2(n1211), .ZN(n1212) );
  CKND0BWP U740 ( .I(n1213), .ZN(n1207) );
  CKND2D0BWP U741 ( .A1(n755), .A2(n1192), .ZN(n1205) );
  CKND2D0BWP U742 ( .A1(n1159), .A2(n1158), .ZN(n1222) );
  CKND2D0BWP U743 ( .A1(n1157), .A2(n1184), .ZN(n1158) );
  CKND0BWP U744 ( .I(n1199), .ZN(n1170) );
  CKND0BWP U745 ( .I(n1152), .ZN(n1155) );
  CKND2D0BWP U746 ( .A1(n1194), .A2(n1192), .ZN(n1196) );
  CKND0BWP U747 ( .I(n1193), .ZN(n1168) );
  CKND2D0BWP U748 ( .A1(n1149), .A2(n1184), .ZN(n1165) );
  CKND2D0BWP U749 ( .A1(n1167), .A2(n1201), .ZN(n1191) );
  CKND0BWP U750 ( .I(n1194), .ZN(n1206) );
  CKND0BWP U751 ( .I(n1184), .ZN(n1164) );
  CKND0BWP U752 ( .I(n1200), .ZN(n755) );
  OR2XD1BWP U753 ( .A1(n1190), .A2(n1208), .Z(n1200) );
  CKND0BWP U754 ( .I(n1161), .ZN(n1156) );
  CKND2D0BWP U755 ( .A1(n1152), .A2(n1154), .ZN(n1162) );
  CKND2D0BWP U756 ( .A1(n1132), .A2(n1149), .ZN(n1147) );
  XOR2D1BWP U757 ( .A1(n1130), .A2(n1136), .Z(n1163) );
  CKND0BWP U758 ( .I(n1132), .ZN(n1151) );
  CKND2D0BWP U759 ( .A1(n1130), .A2(n1181), .ZN(n1123) );
  CKND0BWP U760 ( .I(n1141), .ZN(n1146) );
  CKND0BWP U761 ( .I(n575), .ZN(n564) );
  CKND0BWP U762 ( .I(n1111), .ZN(n1089) );
  CKND0BWP U763 ( .I(n1105), .ZN(n1109) );
  CKND2D0BWP U764 ( .A1(n1104), .A2(n1103), .ZN(n1099) );
  CKND0BWP U765 ( .I(n1102), .ZN(n1128) );
  CKND2D0BWP U766 ( .A1(n1126), .A2(n1122), .ZN(n1124) );
  CKND0BWP U767 ( .I(n1130), .ZN(n1110) );
  CKND2D0BWP U768 ( .A1(n1092), .A2(n1176), .ZN(n1107) );
  MOAI22D0BWP U769 ( .A1(n1120), .A2(n1119), .B1(n1173), .B2(n1177), .ZN(n1121) );
  CKND0BWP U770 ( .I(n1136), .ZN(n1181) );
  CKND2D0BWP U771 ( .A1(n1088), .A2(n1111), .ZN(n1136) );
  CKND0BWP U772 ( .I(n1072), .ZN(n1074) );
  CKND0BWP U773 ( .I(n1071), .ZN(n1101) );
  CKND0BWP U774 ( .I(n1070), .ZN(n1097) );
  CKND0BWP U775 ( .I(n1069), .ZN(n1098) );
  CKND2D0BWP U776 ( .A1(n1062), .A2(n1092), .ZN(n1090) );
  CKND0BWP U777 ( .I(n1095), .ZN(n1106) );
  XOR2D1BWP U778 ( .A1(n1065), .A2(n1173), .Z(n1095) );
  CKND0BWP U779 ( .I(n1062), .ZN(n1094) );
  CKND0BWP U780 ( .I(n1054), .ZN(n1057) );
  CKND0BWP U781 ( .I(n1076), .ZN(n1080) );
  CKND0BWP U782 ( .I(n1042), .ZN(n982) );
  OA222D1BWP U783 ( .A1(n942), .A2(n978), .B1(n941), .B2(n940), .C1(n976), 
        .C2(n1314), .Z(n1043) );
  CKND0BWP U784 ( .I(n1119), .ZN(n1176) );
  OR2XD1BWP U785 ( .A1(n1076), .A2(n1079), .Z(n1119) );
  CKND2D0BWP U786 ( .A1(n1040), .A2(n1039), .ZN(n1076) );
  CKND0BWP U787 ( .I(n1061), .ZN(n1068) );
  CKND0BWP U788 ( .I(n1028), .ZN(n1030) );
  CKND0BWP U789 ( .I(n1027), .ZN(n1031) );
  CKND2D0BWP U790 ( .A1(n1027), .A2(n1028), .ZN(n1023) );
  CKND0BWP U791 ( .I(n1026), .ZN(n1059) );
  CKND2D0BWP U792 ( .A1(n1054), .A2(n1055), .ZN(n1056) );
  XOR2D1BWP U793 ( .A1(n1053), .A2(n1032), .Z(n1065) );
  CKND2D0BWP U794 ( .A1(n1053), .A2(n1017), .ZN(n1033) );
  CKND0BWP U795 ( .I(n1046), .ZN(n979) );
  CKND2D0BWP U796 ( .A1(n1014), .A2(n1040), .ZN(n1173) );
  CKND0BWP U797 ( .I(n997), .ZN(n1022) );
  CKND0BWP U798 ( .I(n996), .ZN(n1021) );
  CKND2D0BWP U799 ( .A1(n758), .A2(n986), .ZN(n992) );
  CKND2D0BWP U800 ( .A1(n983), .A2(n758), .ZN(n985) );
  CKND0BWP U801 ( .I(n1006), .ZN(n628) );
  CKND2D0BWP U802 ( .A1(N115), .A2(n623), .ZN(n624) );
  CKND0BWP U803 ( .I(n691), .ZN(n623) );
  CKND0BWP U804 ( .I(N116), .ZN(n637) );
  CKND2D0BWP U805 ( .A1(n758), .A2(n1116), .ZN(n1118) );
  CKND0BWP U806 ( .I(n1053), .ZN(n1116) );
  CKND2D0BWP U807 ( .A1(n956), .A2(n955), .ZN(n1025) );
  CKND2D0BWP U808 ( .A1(n759), .A2(n954), .ZN(n955) );
  CKND0BWP U809 ( .I(n999), .ZN(n966) );
  CKND0BWP U810 ( .I(n949), .ZN(n951) );
  CKND2D0BWP U811 ( .A1(n986), .A2(n993), .ZN(n990) );
  CKND2D0BWP U812 ( .A1(n963), .A2(n983), .ZN(n984) );
  CKND0BWP U813 ( .I(n988), .ZN(n964) );
  CKND2D0BWP U814 ( .A1(n759), .A2(n946), .ZN(n961) );
  CKND2D0BWP U815 ( .A1(n993), .A2(n994), .ZN(n969) );
  CKND0BWP U816 ( .I(n983), .ZN(n994) );
  CKND0BWP U817 ( .I(n973), .ZN(n975) );
  CKND0BWP U818 ( .I(n640), .ZN(n641) );
  CKND2D0BWP U819 ( .A1(n706), .A2(N1782), .ZN(n640) );
  CKND0BWP U820 ( .I(n757), .ZN(n588) );
  CKND2D0BWP U821 ( .A1(n1051), .A2(n1050), .ZN(n589) );
  CKND0BWP U822 ( .I(n758), .ZN(n1051) );
  CKAN2D0BWP U823 ( .A1(n973), .A2(n974), .Z(n758) );
  CKND0BWP U824 ( .I(N117), .ZN(n713) );
  CKND0BWP U825 ( .I(n939), .ZN(n918) );
  CKND0BWP U826 ( .I(n959), .ZN(n953) );
  CKND0BWP U827 ( .I(n931), .ZN(n933) );
  CKND2D0BWP U828 ( .A1(n949), .A2(n952), .ZN(n958) );
  XNR2D1BWP U829 ( .A1(n927), .A2(n1084), .ZN(n960) );
  CKND2D0BWP U830 ( .A1(n921), .A2(n1319), .ZN(n929) );
  CKND0BWP U831 ( .I(n1084), .ZN(n1319) );
  CKND0BWP U832 ( .I(N114), .ZN(n704) );
  CKND0BWP U833 ( .I(n1050), .ZN(n759) );
  OR2XD1BWP U834 ( .A1(n917), .A2(n939), .Z(n1050) );
  CKND2D0BWP U835 ( .A1(n1317), .A2(n901), .ZN(n903) );
  CKND2D0BWP U836 ( .A1(n930), .A2(n921), .ZN(n926) );
  CKAN2D0BWP U837 ( .A1(n919), .A2(n923), .Z(n921) );
  CKND2D0BWP U838 ( .A1(n1317), .A2(n894), .ZN(n902) );
  CKND0BWP U839 ( .I(n890), .ZN(n892) );
  CKND2D0BWP U840 ( .A1(n766), .A2(n1315), .ZN(n1048) );
  CKND0BWP U841 ( .I(N118), .ZN(n651) );
  CKND0BWP U842 ( .I(n1317), .ZN(n1315) );
  MOAI22D0BWP U843 ( .A1(n940), .A2(n1314), .B1(n912), .B2(n562), .ZN(n558) );
  MAOI22D0BWP U844 ( .A1(n752), .A2(n700), .B1(n597), .B2(N115), .ZN(n556) );
  CKND0BWP U845 ( .I(N113), .ZN(n700) );
  CKND2D0BWP U846 ( .A1(n1317), .A2(n1084), .ZN(n981) );
  MOAI22D0BWP U847 ( .A1(n941), .A2(n697), .B1(n698), .B2(n570), .ZN(n571) );
  CKND0BWP U848 ( .I(N108), .ZN(n682) );
  CKND0BWP U849 ( .I(n699), .ZN(n572) );
  CKND0BWP U850 ( .I(N111), .ZN(n694) );
  CKND0BWP U851 ( .I(N110), .ZN(n688) );
  CKND0BWP U852 ( .I(n597), .ZN(n683) );
  CKND0BWP U853 ( .I(N109), .ZN(n686) );
  CKND0BWP U854 ( .I(n942), .ZN(n912) );
  CKND2D0BWP U855 ( .A1(n1314), .A2(n941), .ZN(n942) );
  CKND2D0BWP U856 ( .A1(n911), .A2(n910), .ZN(n1084) );
  CKND0BWP U857 ( .I(n885), .ZN(n887) );
  CKND0BWP U858 ( .I(N119), .ZN(n657) );
  CKND0BWP U859 ( .I(N123), .ZN(n671) );
  CKND0BWP U860 ( .I(n609), .ZN(n633) );
  CKND0BWP U861 ( .I(N120), .ZN(n662) );
  CKND0BWP U862 ( .I(n632), .ZN(n684) );
  CKND0BWP U863 ( .I(n880), .ZN(n882) );
  CKND0BWP U864 ( .I(n900), .ZN(n897) );
  CKND2D0BWP U865 ( .A1(n890), .A2(n893), .ZN(n900) );
  CKAN2D0BWP U866 ( .A1(n901), .A2(n879), .Z(n894) );
  XOR2D1BWP U867 ( .A1(n876), .A2(n941), .Z(n901) );
  CKND2D0BWP U868 ( .A1(n868), .A2(n766), .ZN(n875) );
  CKND0BWP U869 ( .I(n877), .ZN(n869) );
  CKND2D0BWP U870 ( .A1(n766), .A2(n867), .ZN(n877) );
  CKND2D0BWP U871 ( .A1(n885), .A2(n886), .ZN(n941) );
  CKND0BWP U872 ( .I(N122), .ZN(n669) );
  CKND0BWP U873 ( .I(N121), .ZN(n667) );
  CKND0BWP U874 ( .I(n864), .ZN(n866) );
  CKND2D0BWP U875 ( .A1(n885), .A2(n863), .ZN(n909) );
  CKND0BWP U876 ( .I(n898), .ZN(n860) );
  CKND2D0BWP U877 ( .A1(n874), .A2(n868), .ZN(n873) );
  CKAN2D0BWP U878 ( .A1(n867), .A2(n870), .Z(n868) );
  CKND2D0BWP U879 ( .A1(n1314), .A2(n850), .ZN(n857) );
  XOR2D1BWP U880 ( .A1(n856), .A2(n1314), .Z(n876) );
  CKND0BWP U881 ( .I(n1314), .ZN(n698) );
  CKAN2D0BWP U882 ( .A1(n845), .A2(n1314), .Z(n851) );
  CKND0BWP U883 ( .I(N124), .ZN(n674) );
  CKND2D0BWP U884 ( .A1(n597), .A2(n913), .ZN(n632) );
  CKND2D0BWP U885 ( .A1(n752), .A2(n1313), .ZN(n691) );
  CKND2D0BWP U886 ( .A1(n844), .A2(n840), .ZN(n864) );
  CKND2D0BWP U887 ( .A1(n832), .A2(n831), .ZN(n833) );
  CKND2D0BWP U888 ( .A1(n846), .A2(n856), .ZN(n828) );
  CKND2D0BWP U889 ( .A1(n846), .A2(n845), .ZN(n848) );
  XOR2D1BWP U890 ( .A1(n831), .A2(n762), .Z(n856) );
  XNR2D1BWP U891 ( .A1(n832), .A2(n822), .ZN(n846) );
  MUX2D1BWP U892 ( .I0(n820), .I1(n826), .S(n1313), .Z(n830) );
  CKND2D0BWP U893 ( .A1(n832), .A2(n819), .ZN(n829) );
  CKND2D0BWP U894 ( .A1(n819), .A2(n762), .ZN(n822) );
  CKND0BWP U895 ( .I(n814), .ZN(n839) );
  CKND0BWP U896 ( .I(n816), .ZN(n809) );
  CKND0BWP U897 ( .I(n762), .ZN(n1009) );
  CKAN2D0BWP U898 ( .A1(n763), .A2(n844), .Z(n762) );
  CKND2D0BWP U899 ( .A1(n794), .A2(n752), .ZN(n796) );
  CKND0BWP U900 ( .I(n800), .ZN(n793) );
  CKND2D0BWP U901 ( .A1(n795), .A2(n794), .ZN(n801) );
  CKND0BWP U902 ( .I(n823), .ZN(n837) );
  CKND2D0BWP U903 ( .A1(n761), .A2(n799), .ZN(n812) );
  CKND2D0BWP U904 ( .A1(n761), .A2(n807), .ZN(n791) );
  CKND2D0BWP U905 ( .A1(n599), .A2(n598), .ZN(n602) );
  CKND0BWP U906 ( .I(n786), .ZN(n598) );
  XNR2D1BWP U907 ( .A1(n599), .A2(n786), .ZN(n795) );
  CKND0BWP U908 ( .I(n788), .ZN(n798) );
  CKND2D0BWP U909 ( .A1(n789), .A2(n783), .ZN(n787) );
  CKND2D0BWP U910 ( .A1(n752), .A2(n789), .ZN(n784) );
  CKND0BWP U911 ( .I(n913), .ZN(n752) );
  CKND0BWP U912 ( .I(n1238), .ZN(n642) );
  CKND2D0BWP U913 ( .A1(n1238), .A2(n780), .ZN(n777) );
  CKND2D0BWP U914 ( .A1(n774), .A2(n709), .ZN(n548) );
  CKND0BWP U915 ( .I(n1344), .ZN(n1341) );
  CKND0BWP U916 ( .I(n1343), .ZN(n1308) );
  CKND2D0BWP U917 ( .A1(n593), .A2(n594), .ZN(n783) );
  CKND2D0BWP U918 ( .A1(n597), .A2(n595), .ZN(n594) );
  CKND0BWP U919 ( .I(n592), .ZN(n595) );
  CKND2D0BWP U920 ( .A1(n774), .A2(n1334), .ZN(n778) );
  CKND0BWP U921 ( .I(n1333), .ZN(n1334) );
  CKND2D0BWP U922 ( .A1(n709), .A2(n708), .ZN(n549) );
  CKND0BWP U923 ( .I(N126), .ZN(n708) );
  CKND0BWP U924 ( .I(n596), .ZN(n593) );
  CKND0BWP U925 ( .I(n1335), .ZN(n1328) );
  CKND0BWP U926 ( .I(N1940), .ZN(n646) );
  CKND0BWP U927 ( .I(N127), .ZN(n709) );
  CKND2D0BWP U928 ( .A1(A[13]), .A2(n1322), .ZN(n1349) );
  AN4D1BWP U929 ( .A1(A[10]), .A2(A[11]), .A3(A[14]), .A4(A[12]), .Z(n1322) );
  CKND2D0BWP U930 ( .A1(n639), .A2(n655), .ZN(n1324) );
  CKND2D0BWP U931 ( .A1(N1940), .A2(n1323), .ZN(n655) );
  CKND0BWP U932 ( .I(A[1]), .ZN(n537) );
  CKND0BWP U933 ( .I(A[3]), .ZN(n538) );
  CKND0BWP U934 ( .I(A[5]), .ZN(n539) );
  CKND0BWP U935 ( .I(\DP_OP_379J1_125_371/n49 ), .ZN(n545) );
  CKND0BWP U936 ( .I(A[9]), .ZN(n541) );
  CKND0BWP U937 ( .I(B[8]), .ZN(n533) );
  CKND0BWP U938 ( .I(N93), .ZN(n535) );
  CKND0BWP U939 ( .I(n1325), .ZN(n639) );
  CKND2D0BWP U940 ( .A1(n1344), .A2(n1343), .ZN(n1239) );
  CKND2D0BWP U941 ( .A1(n1333), .A2(n1335), .ZN(n1338) );
  CKND2D0BWP U942 ( .A1(n765), .A2(n767), .ZN(n768) );
  XNR2D1BWP U943 ( .A1(n755), .A2(n1201), .ZN(n1223) );
  XNR2D1BWP U944 ( .A1(n1184), .A2(n1163), .ZN(n1201) );
  XNR2D1BWP U945 ( .A1(n1317), .A2(n901), .ZN(n927) );
  XNR2D1BWP U946 ( .A1(n1256), .A2(n1251), .ZN(n1270) );
  NR3D0BWP U947 ( .A1(n1325), .A2(N78), .A3(n655), .ZN(n749) );
  NR2XD0BWP U948 ( .A1(n649), .A2(n741), .ZN(\DP_OP_379J1_125_371/I5 ) );
  NR2XD0BWP U949 ( .A1(n1141), .A2(n1145), .ZN(n1184) );
  XNR2D1BWP U950 ( .A1(n1064), .A2(n1063), .ZN(n1091) );
  XNR2D1BWP U951 ( .A1(n1016), .A2(n1018), .ZN(n1064) );
  NR2XD0BWP U952 ( .A1(n746), .A2(n641), .ZN(n712) );
  MOAI22D0BWP U953 ( .A1(n940), .A2(n942), .B1(n766), .B2(n562), .ZN(n563) );
  XNR2D1BWP U954 ( .A1(n889), .A2(n895), .ZN(n930) );
  NR2XD0BWP U955 ( .A1(n909), .A2(n908), .ZN(n1317) );
  NR2XD0BWP U956 ( .A1(n864), .A2(n865), .ZN(n1314) );
  NR2XD0BWP U957 ( .A1(n549), .A2(n782), .ZN(n597) );
  ND2D1BWP U958 ( .A1(n709), .A2(n646), .ZN(n746) );
  NR2XD0BWP U959 ( .A1(n1324), .A2(N78), .ZN(n750) );
  AOI21D1BWP U960 ( .A1(n776), .A2(B[14]), .B(n1310), .ZN(n1238) );
  FA1D0BWP U961 ( .A(A[13]), .B(B[13]), .CI(n770), .CO(n771), .S(n1344) );
  NR2XD0BWP U962 ( .A1(n722), .A2(n721), .ZN(n745) );
  NR2XD0BWP U963 ( .A1(n1241), .A2(n1240), .ZN(n756) );
  NR2XD0BWP U964 ( .A1(n1004), .A2(n1005), .ZN(n1053) );
  OAI31D1BWP U965 ( .A1(n969), .A2(n968), .A3(n967), .B(n973), .ZN(n1005) );
  AOI31D1BWP U966 ( .A1(n820), .A2(n805), .A3(n824), .B(n806), .ZN(n844) );
  INVD1BWP U967 ( .I(B[14]), .ZN(n764) );
  INVD1BWP U968 ( .I(n1326), .ZN(n1337) );
  OAI21D1BWP U969 ( .A1(n767), .A2(n765), .B(n768), .ZN(n1326) );
  INVD1BWP U970 ( .I(A[10]), .ZN(n767) );
  IND2D1BWP U971 ( .A1(N78), .B1(n1324), .ZN(N1942) );
  OAI31D1BWP U972 ( .A1(n1318), .A2(n1319), .A3(n546), .B(n705), .ZN(N1927) );
  AOI22D1BWP U973 ( .A1(n1317), .A2(n760), .B1(n1316), .B2(n1315), .ZN(n1318)
         );
  MUX2ND0BWP U974 ( .I0(n682), .I1(n681), .S(n751), .ZN(N1920) );
  MUX2D1BWP U975 ( .I0(N124), .I1(N1789), .S(n751), .Z(N1936) );
  MUX2ND0BWP U976 ( .I0(n708), .I1(n707), .S(n751), .ZN(N1938) );
  OAI21D1BWP U977 ( .A1(n1312), .A2(n546), .B(n1311), .ZN(N1917) );
  AO21D1BWP U978 ( .A1(n751), .A2(n1309), .B(n642), .Z(N1916) );
  AOI22D1BWP U979 ( .A1(n751), .A2(n1345), .B1(n1308), .B2(n546), .ZN(N1915)
         );
  OAI21D1BWP U980 ( .A1(n751), .A2(n704), .B(n703), .ZN(N1926) );
  ND3D1BWP U981 ( .A1(n751), .A2(n760), .A3(n1315), .ZN(n703) );
  AOI22D1BWP U982 ( .A1(n751), .A2(n1342), .B1(n1341), .B2(n546), .ZN(N1914)
         );
  MUX2D1BWP U983 ( .I0(N119), .I1(N1784), .S(n751), .Z(N1931) );
  AOI32D1BWP U984 ( .A1(n1332), .A2(n751), .A3(n1331), .B1(n1334), .B2(n546), 
        .ZN(N1913) );
  MUX2D1BWP U985 ( .I0(N118), .I1(N1783), .S(n751), .Z(N1930) );
  AOI22D1BWP U986 ( .A1(n751), .A2(n1330), .B1(n1328), .B2(n546), .ZN(N1912)
         );
  MUX2D1BWP U987 ( .I0(N117), .I1(N1782), .S(n751), .Z(N1929) );
  AOI22D1BWP U988 ( .A1(n751), .A2(n1327), .B1(n1337), .B2(n546), .ZN(N1911)
         );
  MUX2D1BWP U989 ( .I0(N116), .I1(n706), .S(n751), .Z(N1928) );
  MUX2D1BWP U990 ( .I0(N123), .I1(N1788), .S(n751), .Z(N1935) );
  MUX2D1BWP U991 ( .I0(N122), .I1(N1787), .S(n751), .Z(N1934) );
  MUX2D1BWP U992 ( .I0(N121), .I1(N1786), .S(n751), .Z(N1933) );
  OAI22D1BWP U993 ( .A1(n702), .A2(n701), .B1(n751), .B2(n700), .ZN(N1925) );
  AOI22D1BWP U994 ( .A1(n699), .A2(n698), .B1(n697), .B2(n1314), .ZN(n702) );
  MUX2D1BWP U995 ( .I0(N120), .I1(N1785), .S(n751), .Z(N1932) );
  OAI31D1BWP U996 ( .A1(n1314), .A2(n546), .A3(n696), .B(n695), .ZN(N1924) );
  OAI22D1BWP U997 ( .A1(n751), .A2(n694), .B1(n693), .B2(n692), .ZN(N1923) );
  OAI22D1BWP U998 ( .A1(N108), .A2(n691), .B1(n690), .B2(n1313), .ZN(n692) );
  OAI211D1BWP U999 ( .A1(n761), .A2(n689), .B(n751), .C(n1009), .ZN(n693) );
  OAI21D1BWP U1000 ( .A1(n1320), .A2(n546), .B(n709), .ZN(N1939) );
  OAI21D1BWP U1001 ( .A1(n751), .A2(n688), .B(n687), .ZN(N1922) );
  ND3D1BWP U1002 ( .A1(n751), .A2(n690), .A3(n1313), .ZN(n687) );
  MUX2ND0BWP U1003 ( .I0(n686), .I1(n685), .S(n751), .ZN(N1921) );
  AOI22D1BWP U1004 ( .A1(N107), .A2(n684), .B1(N108), .B2(n683), .ZN(n685) );
  MUX2D1BWP U1005 ( .I0(N125), .I1(N1790), .S(n751), .Z(N1937) );
  OAI221D1BWP U1006 ( .A1(n1350), .A2(n1349), .B1(n1348), .B2(B[15]), .C(n1347), .ZN(prod[15]) );
  ND3D1BWP U1007 ( .A1(B[15]), .A2(n1349), .A3(n1348), .ZN(n1347) );
  AO22D1BWP U1008 ( .A1(n750), .A2(N1846), .B1(n749), .B2(operprod1[0]), .Z(
        prod[0]) );
  AO21D1BWP U1009 ( .A1(\C148/DATA4_0 ), .A2(n719), .B(n718), .Z(N1846) );
  ND4D1BWP U1010 ( .A1(n717), .A2(n716), .A3(n715), .A4(n720), .ZN(n718) );
  OAI211D1BWP U1011 ( .A1(n651), .A2(n713), .B(N118), .C(n731), .ZN(n715) );
  AO22D1BWP U1012 ( .A1(n750), .A2(N1848), .B1(n749), .B2(operprod1[2]), .Z(
        prod[2]) );
  IOA21D1BWP U1013 ( .A1(\C148/DATA4_2 ), .A2(n719), .B(n660), .ZN(N1848) );
  AOI211XD0BWP U1014 ( .A1(N1784), .A2(n712), .B(n659), .C(n658), .ZN(n660) );
  OAI22D1BWP U1015 ( .A1(n661), .A2(n736), .B1(n673), .B2(n657), .ZN(n658) );
  NR2XD0BWP U1016 ( .A1(n735), .A2(n656), .ZN(n659) );
  AO22D1BWP U1017 ( .A1(n750), .A2(N1849), .B1(n749), .B2(operprod1[3]), .Z(
        prod[3]) );
  IOA21D1BWP U1018 ( .A1(n712), .A2(N1785), .B(n665), .ZN(N1849) );
  AOI211XD0BWP U1019 ( .A1(\C148/DATA4_3 ), .A2(n719), .B(n664), .C(n663), 
        .ZN(n665) );
  OAI22D1BWP U1020 ( .A1(n666), .A2(n736), .B1(n673), .B2(n662), .ZN(n663) );
  NR2XD0BWP U1021 ( .A1(n735), .A2(n661), .ZN(n664) );
  MUX2ND0BWP U1022 ( .I0(N121), .I1(N143), .S(n675), .ZN(n661) );
  AO22D1BWP U1023 ( .A1(n750), .A2(N1850), .B1(n749), .B2(operprod1[4]), .Z(
        prod[4]) );
  MUX2ND0BWP U1024 ( .I0(N122), .I1(N144), .S(n675), .ZN(n666) );
  AO22D1BWP U1025 ( .A1(n750), .A2(N1851), .B1(n749), .B2(operprod1[5]), .Z(
        prod[5]) );
  MUX2ND0BWP U1026 ( .I0(N123), .I1(N145), .S(n675), .ZN(n668) );
  AO22D1BWP U1027 ( .A1(n750), .A2(N1852), .B1(n749), .B2(operprod1[6]), .Z(
        prod[6]) );
  MUX2ND0BWP U1028 ( .I0(N124), .I1(N146), .S(n675), .ZN(n670) );
  AO22D1BWP U1029 ( .A1(n750), .A2(N1853), .B1(n749), .B2(operprod1[7]), .Z(
        prod[7]) );
  MUX2ND0BWP U1030 ( .I0(N125), .I1(N147), .S(n675), .ZN(n672) );
  AO22D1BWP U1031 ( .A1(n750), .A2(N1847), .B1(n749), .B2(operprod1[1]), .Z(
        prod[1]) );
  IOA21D1BWP U1032 ( .A1(\C148/DATA4_1 ), .A2(n719), .B(n654), .ZN(N1847) );
  AOI211XD0BWP U1033 ( .A1(N1783), .A2(n712), .B(n653), .C(n652), .ZN(n654) );
  OAI22D1BWP U1034 ( .A1(n656), .A2(n736), .B1(n651), .B2(n673), .ZN(n652) );
  MUX2ND0BWP U1035 ( .I0(N120), .I1(N142), .S(n675), .ZN(n656) );
  NR2XD0BWP U1036 ( .A1(n735), .A2(n710), .ZN(n653) );
  MUX2ND0BWP U1037 ( .I0(N141), .I1(N119), .S(n647), .ZN(n710) );
  AO22D1BWP U1038 ( .A1(n750), .A2(N1855), .B1(n749), .B2(operprod1[9]), .Z(
        prod[9]) );
  OAI211D1BWP U1039 ( .A1(n1327), .A2(n746), .B(n745), .C(n724), .ZN(prod[10])
         );
  OAI22D1BWP U1040 ( .A1(n730), .A2(n723), .B1(n1326), .B2(n731), .ZN(n724) );
  AOI211XD0BWP U1041 ( .A1(n1306), .A2(n1305), .B(n1304), .C(n1303), .ZN(n1327) );
  IND4D1BWP U1042 ( .A1(n1320), .B1(n1312), .B2(n1345), .B3(n1331), .ZN(n1302)
         );
  IOA21D1BWP U1043 ( .A1(n1298), .A2(n1297), .B(n1296), .ZN(n1309) );
  OAI31D1BWP U1044 ( .A1(n1295), .A2(n1294), .A3(n1293), .B(n1292), .ZN(n1296)
         );
  OAI21D1BWP U1045 ( .A1(n1295), .A2(n1293), .B(n1294), .ZN(n1292) );
  AOI211XD0BWP U1046 ( .A1(n731), .A2(n1329), .B(n726), .C(n725), .ZN(n727) );
  AOI22D1BWP U1047 ( .A1(n1328), .A2(n736), .B1(n1335), .B2(n741), .ZN(n725)
         );
  NR2XD0BWP U1048 ( .A1(n746), .A2(n1330), .ZN(n726) );
  OAI31D1BWP U1049 ( .A1(n1281), .A2(n1303), .A3(n1280), .B(n1279), .ZN(n1330)
         );
  MAOI222D1BWP U1050 ( .A(n1281), .B(n1303), .C(n1280), .ZN(n1279) );
  AO21D1BWP U1051 ( .A1(n1333), .A2(n734), .B(n733), .Z(prod[12]) );
  OAI211D1BWP U1052 ( .A1(n1336), .A2(n746), .B(n745), .C(n732), .ZN(n733) );
  IND3D1BWP U1053 ( .A1(n737), .B1(n1334), .B2(n1335), .ZN(n732) );
  OAI211D1BWP U1054 ( .A1(n729), .A2(n1335), .B(n741), .C(n728), .ZN(n734) );
  OAI211D1BWP U1055 ( .A1(n1342), .A2(n746), .B(n745), .C(n740), .ZN(prod[13])
         );
  OAI22D1BWP U1056 ( .A1(n739), .A2(n738), .B1(n1344), .B2(n748), .ZN(n740) );
  OAI211D1BWP U1057 ( .A1(n1340), .A2(n736), .B(n741), .C(n1344), .ZN(n738) );
  NR2XD0BWP U1058 ( .A1(n735), .A2(n1339), .ZN(n739) );
  NR2XD0BWP U1059 ( .A1(n1338), .A2(n1337), .ZN(n1339) );
  AOI21D1BWP U1060 ( .A1(n1297), .A2(n1290), .B(n1289), .ZN(n1307) );
  OAI21D1BWP U1061 ( .A1(n1297), .A2(n1290), .B(n1332), .ZN(n1289) );
  NR2XD0BWP U1062 ( .A1(n1288), .A2(n1287), .ZN(n1300) );
  AOI31D1BWP U1063 ( .A1(n1298), .A2(n1312), .A3(n1277), .B(n1305), .ZN(n1278)
         );
  OA21D1BWP U1064 ( .A1(n1269), .A2(n756), .B(n1268), .Z(n1312) );
  NR2XD0BWP U1065 ( .A1(n1290), .A2(n1299), .ZN(n1298) );
  AOI21D1BWP U1066 ( .A1(n1272), .A2(n1282), .B(n1275), .ZN(n1286) );
  XOR2D1BWP U1067 ( .A1(n1284), .A2(n1283), .Z(n1301) );
  XOR2D1BWP U1068 ( .A1(n1264), .A2(n1274), .Z(n1290) );
  NR2XD0BWP U1069 ( .A1(n1283), .A2(n1284), .ZN(n1297) );
  OAI21D1BWP U1070 ( .A1(n1276), .A2(n1275), .B(n1274), .ZN(n1284) );
  NR2XD0BWP U1071 ( .A1(n1271), .A2(n1295), .ZN(n1275) );
  IND2D1BWP U1072 ( .A1(n1282), .B1(n1281), .ZN(n1283) );
  NR2XD0BWP U1073 ( .A1(n1305), .A2(n1306), .ZN(n1281) );
  XNR2D1BWP U1074 ( .A1(n756), .A2(n1270), .ZN(n1306) );
  OAI31D1BWP U1075 ( .A1(n1258), .A2(n1257), .A3(n1256), .B(n1255), .ZN(n1261)
         );
  OAI21D1BWP U1076 ( .A1(n1258), .A2(n1256), .B(n1257), .ZN(n1255) );
  NR2XD0BWP U1077 ( .A1(n1266), .A2(n1267), .ZN(n1291) );
  AOI21D1BWP U1078 ( .A1(n1262), .A2(n638), .B(n1241), .ZN(n1320) );
  MUX2ND0BWP U1079 ( .I0(n1234), .I1(n578), .S(n1250), .ZN(n638) );
  XNR2D1BWP U1080 ( .A1(n1260), .A2(n1259), .ZN(n1282) );
  AO21D1BWP U1081 ( .A1(n1344), .A2(n748), .B(n747), .Z(prod[14]) );
  OAI211D1BWP U1082 ( .A1(n1345), .A2(n746), .B(n745), .C(n744), .ZN(n747) );
  OAI21D1BWP U1083 ( .A1(n743), .A2(n742), .B(n1343), .ZN(n744) );
  OAI31D1BWP U1084 ( .A1(n1266), .A2(n1267), .A3(n1295), .B(n1265), .ZN(n1299)
         );
  OAI21D1BWP U1085 ( .A1(n1295), .A2(n1266), .B(n1267), .ZN(n1265) );
  OAI31D1BWP U1086 ( .A1(n1231), .A2(n1230), .A3(n1229), .B(n1228), .ZN(n1254)
         );
  OAI21D1BWP U1087 ( .A1(n1231), .A2(n1229), .B(n1230), .ZN(n1228) );
  IAO21D1BWP U1088 ( .A1(n1222), .A2(n1221), .B(n1220), .ZN(n1269) );
  OAI21D1BWP U1089 ( .A1(n1235), .A2(n1234), .B(n1233), .ZN(n1241) );
  MUX2ND0BWP U1090 ( .I0(n1210), .I1(n577), .S(n1221), .ZN(n1234) );
  OA31D1BWP U1091 ( .A1(n1245), .A2(n1244), .A3(n1256), .B(n1243), .Z(n1267)
         );
  OAI21D1BWP U1092 ( .A1(n1245), .A2(n1256), .B(n1244), .ZN(n1243) );
  OAI31D1BWP U1093 ( .A1(n1216), .A2(n1215), .A3(n1229), .B(n1214), .ZN(n1244)
         );
  OAI21D1BWP U1094 ( .A1(n1216), .A2(n1229), .B(n1215), .ZN(n1214) );
  NR2XD0BWP U1095 ( .A1(n1249), .A2(n1246), .ZN(n1242) );
  NR2XD0BWP U1096 ( .A1(n1271), .A2(n1273), .ZN(n1263) );
  OAI21D1BWP U1097 ( .A1(n1226), .A2(n1225), .B(n1224), .ZN(n1260) );
  NR2XD0BWP U1098 ( .A1(n1229), .A2(n1223), .ZN(n1225) );
  OAI31D1BWP U1099 ( .A1(n1249), .A2(n1248), .A3(n1256), .B(n1247), .ZN(n1264)
         );
  OAI21D1BWP U1100 ( .A1(n1249), .A2(n1256), .B(n1248), .ZN(n1247) );
  XNR2D1BWP U1101 ( .A1(n1219), .A2(n1218), .ZN(n1246) );
  XOR2D1BWP U1102 ( .A1(n1223), .A2(n1229), .Z(n1251) );
  AOI21D1BWP U1103 ( .A1(n1213), .A2(n1224), .B(n1218), .ZN(n1252) );
  NR2XD0BWP U1104 ( .A1(n1229), .A2(n1212), .ZN(n1218) );
  NR2XD0BWP U1105 ( .A1(n1338), .A2(n737), .ZN(n748) );
  AOI21D1BWP U1106 ( .A1(n731), .A2(n1326), .B(n730), .ZN(n737) );
  AO22D1BWP U1107 ( .A1(n750), .A2(N1854), .B1(n749), .B2(operprod1[8]), .Z(
        prod[8]) );
  AO21D1BWP U1108 ( .A1(n712), .A2(N1790), .B(n679), .Z(N1854) );
  OAI211D1BWP U1109 ( .A1(n678), .A2(n735), .B(n677), .C(n676), .ZN(n679) );
  OR2XD1BWP U1110 ( .A1(\DP_OP_379J1_125_371/I4 ), .A2(
        \DP_OP_379J1_125_371/I5 ), .Z(n719) );
  AOI211XD0BWP U1111 ( .A1(n1119), .A2(n584), .B(n583), .C(n1181), .ZN(N1786)
         );
  NR2XD0BWP U1112 ( .A1(n1119), .A2(n585), .ZN(n583) );
  NR2XD0BWP U1113 ( .A1(n582), .A2(n1184), .ZN(N1787) );
  AOI211XD0BWP U1114 ( .A1(n1184), .A2(n582), .B(n755), .C(n581), .ZN(N1788)
         );
  NR2XD0BWP U1115 ( .A1(n580), .A2(n1184), .ZN(n581) );
  NR2XD0BWP U1116 ( .A1(n640), .A2(n746), .ZN(\DP_OP_379J1_125_371/I4 ) );
  MUX2ND0BWP U1117 ( .I0(N127), .I1(N149), .S(n675), .ZN(n680) );
  NR2XD0BWP U1118 ( .A1(n741), .A2(n650), .ZN(n711) );
  NR3D0BWP U1119 ( .A1(n714), .A2(n648), .A3(n646), .ZN(n731) );
  NR4D0BWP U1120 ( .A1(n1237), .A2(n1323), .A3(n647), .A4(n645), .ZN(n648) );
  AOI21D1BWP U1121 ( .A1(n644), .A2(n643), .B(n642), .ZN(n714) );
  ND4D1BWP U1122 ( .A1(n675), .A2(n1237), .A3(\DP_OP_379J1_125_371/n10 ), .A4(
        n1328), .ZN(n643) );
  OAI211D1BWP U1123 ( .A1(N150), .A2(n647), .B(n1337), .C(n1236), .ZN(n644) );
  NR2XD0BWP U1124 ( .A1(n1239), .A2(n1338), .ZN(n1236) );
  MUX2ND0BWP U1125 ( .I0(N126), .I1(N148), .S(n675), .ZN(n678) );
  NR2XD0BWP U1126 ( .A1(n578), .A2(n1250), .ZN(N1790) );
  NR2XD0BWP U1127 ( .A1(n1190), .A2(n1189), .ZN(n1233) );
  OAI32D1BWP U1128 ( .A1(n1208), .A2(n1209), .A3(n1188), .B1(n754), .B2(n1208), 
        .ZN(n1189) );
  AOI21D1BWP U1129 ( .A1(n1204), .A2(n1203), .B(n1202), .ZN(n1226) );
  IND2D1BWP U1130 ( .A1(n1216), .B1(n1215), .ZN(n1231) );
  OAI31D1BWP U1131 ( .A1(n1200), .A2(n1197), .A3(n1196), .B(n1195), .ZN(n1215)
         );
  OAI21D1BWP U1132 ( .A1(n1200), .A2(n1196), .B(n1197), .ZN(n1195) );
  IND2D1BWP U1133 ( .A1(n1212), .B1(n1219), .ZN(n1216) );
  NR2XD0BWP U1134 ( .A1(n1203), .A2(n1223), .ZN(n1211) );
  OAI21D1BWP U1135 ( .A1(n1193), .A2(n1202), .B(n1205), .ZN(n1213) );
  NR2XD0BWP U1136 ( .A1(n1191), .A2(n1200), .ZN(n1202) );
  MUX2ND0BWP U1137 ( .I0(n577), .I1(n579), .S(n1221), .ZN(n578) );
  INR3D0BWP U1138 ( .A1(n754), .B1(n1209), .B2(n1200), .ZN(n1221) );
  OAI211D1BWP U1139 ( .A1(n1170), .A2(n1222), .B(n1198), .C(n1169), .ZN(n1171)
         );
  AOI21D1BWP U1140 ( .A1(n1168), .A2(n1191), .B(n1203), .ZN(n1169) );
  OAI21D1BWP U1141 ( .A1(n1167), .A2(n1166), .B(n1165), .ZN(n1203) );
  NR2XD0BWP U1142 ( .A1(n1164), .A2(n1163), .ZN(n1166) );
  OAI31D1BWP U1143 ( .A1(n1162), .A2(n1161), .A3(n1164), .B(n1160), .ZN(n1198)
         );
  OAI21D1BWP U1144 ( .A1(n1162), .A2(n1164), .B(n1161), .ZN(n1160) );
  NR2XD0BWP U1145 ( .A1(n1162), .A2(n1156), .ZN(n1157) );
  IND2D1BWP U1146 ( .A1(n1196), .B1(n1197), .ZN(n1199) );
  XOR2D1BWP U1147 ( .A1(n1196), .A2(n1197), .Z(n1172) );
  OAI31D1BWP U1148 ( .A1(n1155), .A2(n1154), .A3(n1164), .B(n1153), .ZN(n1197)
         );
  OAI21D1BWP U1149 ( .A1(n1155), .A2(n1164), .B(n1154), .ZN(n1153) );
  NR2XD0BWP U1150 ( .A1(n1191), .A2(n1168), .ZN(n1192) );
  AOI21D1BWP U1151 ( .A1(n1151), .A2(n1165), .B(n1150), .ZN(n1193) );
  XNR2D1BWP U1152 ( .A1(n1148), .A2(n1150), .ZN(n1194) );
  NR2XD0BWP U1153 ( .A1(n1164), .A2(n1147), .ZN(n1150) );
  MUX2ND0BWP U1154 ( .I0(n1180), .I1(n1186), .S(n1184), .ZN(n754) );
  MUX2ND0BWP U1155 ( .I0(n576), .I1(n582), .S(n755), .ZN(n579) );
  MUX2ND0BWP U1156 ( .I0(n575), .I1(n585), .S(n1181), .ZN(n582) );
  MUX2ND0BWP U1157 ( .I0(n574), .I1(n573), .S(n1053), .ZN(n585) );
  MUX2ND0BWP U1158 ( .I0(n587), .I1(n586), .S(n1173), .ZN(n573) );
  AOI222D1BWP U1159 ( .A1(n591), .A2(n758), .B1(n590), .B2(n757), .C1(n1050), 
        .C2(n1044), .ZN(n587) );
  MUX2ND0BWP U1160 ( .I0(n1187), .I1(n576), .S(n755), .ZN(n577) );
  IND2D1BWP U1161 ( .A1(n1142), .B1(n1146), .ZN(n1208) );
  AO211D1BWP U1162 ( .A1(n1162), .A2(n1159), .B(n1156), .C(n1138), .Z(n1139)
         );
  IND2D1BWP U1163 ( .A1(n1148), .B1(n1163), .ZN(n1138) );
  XNR2D1BWP U1164 ( .A1(n1154), .A2(n1152), .ZN(n1140) );
  NR2XD0BWP U1165 ( .A1(n1147), .A2(n1148), .ZN(n1152) );
  XNR2D1BWP U1166 ( .A1(n1134), .A2(n1133), .ZN(n1148) );
  NR2XD0BWP U1167 ( .A1(n1163), .A2(n1131), .ZN(n1149) );
  OAI31D1BWP U1168 ( .A1(n1129), .A2(n1128), .A3(n1136), .B(n1127), .ZN(n1154)
         );
  OAI21D1BWP U1169 ( .A1(n1129), .A2(n1136), .B(n1128), .ZN(n1127) );
  IAO21D1BWP U1170 ( .A1(n1126), .A2(n1125), .B(n1133), .ZN(n1132) );
  NR2XD0BWP U1171 ( .A1(n1124), .A2(n1136), .ZN(n1133) );
  AOI21D1BWP U1172 ( .A1(n1131), .A2(n1123), .B(n1125), .ZN(n1167) );
  INR2D1BWP U1173 ( .A1(n1122), .B1(n1136), .ZN(n1125) );
  AO21D1BWP U1174 ( .A1(n1146), .A2(n1180), .B(n1145), .Z(n1190) );
  MUX2ND0BWP U1175 ( .I0(n1185), .I1(n580), .S(n1184), .ZN(n576) );
  MUX2ND0BWP U1176 ( .I0(n1182), .I1(n564), .S(n1181), .ZN(n580) );
  MUX2ND0BWP U1177 ( .I0(n1120), .I1(n584), .S(n1176), .ZN(n575) );
  MUX2D1BWP U1178 ( .I0(n1112), .I1(n574), .S(n1053), .Z(n584) );
  MUX2ND0BWP U1179 ( .I0(n586), .I1(n1113), .S(n1173), .ZN(n574) );
  AOI222D1BWP U1180 ( .A1(n590), .A2(n758), .B1(n757), .B2(n1044), .C1(n1050), 
        .C2(n1052), .ZN(n586) );
  OAI21D1BWP U1181 ( .A1(n1144), .A2(n1089), .B(n1088), .ZN(n1145) );
  AOI222D1BWP U1182 ( .A1(n1087), .A2(n1173), .B1(n1143), .B2(n1178), .C1(
        n1174), .C2(n1176), .ZN(n1144) );
  OAI21D1BWP U1183 ( .A1(n1109), .A2(n1108), .B(n1107), .ZN(n1131) );
  NR2XD0BWP U1184 ( .A1(n1119), .A2(n1106), .ZN(n1108) );
  OR2XD1BWP U1185 ( .A1(n1129), .A2(n1102), .Z(n1137) );
  NR2XD0BWP U1186 ( .A1(n1101), .A2(n1100), .ZN(n1159) );
  NR2XD0BWP U1187 ( .A1(n1119), .A2(n1099), .ZN(n1100) );
  OAI31D1BWP U1188 ( .A1(n1098), .A2(n1097), .A3(n1119), .B(n1096), .ZN(n1102)
         );
  OAI21D1BWP U1189 ( .A1(n1098), .A2(n1119), .B(n1097), .ZN(n1096) );
  IND2D1BWP U1190 ( .A1(n1124), .B1(n1134), .ZN(n1129) );
  NR2XD0BWP U1191 ( .A1(n1105), .A2(n1110), .ZN(n1122) );
  XNR2D1BWP U1192 ( .A1(n1095), .A2(n1119), .ZN(n1130) );
  AOI21D1BWP U1193 ( .A1(n1094), .A2(n1107), .B(n1093), .ZN(n1126) );
  XNR2D1BWP U1194 ( .A1(n1091), .A2(n1093), .ZN(n1134) );
  NR2XD0BWP U1195 ( .A1(n1119), .A2(n1090), .ZN(n1093) );
  AOI21D1BWP U1196 ( .A1(n1178), .A2(n1175), .B(n1121), .ZN(n1182) );
  AOI222D1BWP U1197 ( .A1(n1049), .A2(n1050), .B1(n1052), .B2(n757), .C1(n1044), .C2(n758), .ZN(n1113) );
  OAI222D1BWP U1198 ( .A1(n981), .A2(n980), .B1(n1084), .B2(n943), .C1(n1043), 
        .C2(n1317), .ZN(n1044) );
  OAI31D1BWP U1199 ( .A1(n1075), .A2(n1074), .A3(n1173), .B(n1073), .ZN(n1104)
         );
  OAI21D1BWP U1200 ( .A1(n1075), .A2(n1173), .B(n1074), .ZN(n1073) );
  NR2XD0BWP U1201 ( .A1(n1098), .A2(n1097), .ZN(n1103) );
  OAI21D1BWP U1202 ( .A1(n1068), .A2(n1067), .B(n1066), .ZN(n1105) );
  NR2XD0BWP U1203 ( .A1(n1173), .A2(n1065), .ZN(n1067) );
  NR2XD0BWP U1204 ( .A1(n1090), .A2(n1091), .ZN(n1069) );
  NR2XD0BWP U1205 ( .A1(n1106), .A2(n1061), .ZN(n1092) );
  OAI31D1BWP U1206 ( .A1(n1060), .A2(n1059), .A3(n1173), .B(n1058), .ZN(n1070)
         );
  OAI21D1BWP U1207 ( .A1(n1060), .A2(n1173), .B(n1059), .ZN(n1058) );
  AOI21D1BWP U1208 ( .A1(n1057), .A2(n1066), .B(n1063), .ZN(n1062) );
  NR2XD0BWP U1209 ( .A1(n1056), .A2(n1173), .ZN(n1063) );
  IND2D1BWP U1210 ( .A1(n1173), .B1(n1055), .ZN(n1066) );
  AOI21D1BWP U1211 ( .A1(n1080), .A2(n1143), .B(n1079), .ZN(n1088) );
  AOI222D1BWP U1212 ( .A1(n1178), .A2(n1177), .B1(n1176), .B2(n1175), .C1(
        n1174), .C2(n1173), .ZN(n1183) );
  MUX2D1BWP U1213 ( .I0(n1052), .I1(n1115), .S(n1051), .Z(n1112) );
  OAI222D1BWP U1214 ( .A1(n982), .A2(n1317), .B1(n1043), .B2(n981), .C1(n980), 
        .C2(n1084), .ZN(n1052) );
  AOI222D1BWP U1215 ( .A1(n1143), .A2(n1173), .B1(n1174), .B2(n1178), .C1(
        n1177), .C2(n1176), .ZN(n1179) );
  OAI222D1BWP U1216 ( .A1(n1118), .A2(n1117), .B1(n1116), .B2(n1115), .C1(
        n1114), .C2(n758), .ZN(n1177) );
  NR2XD0BWP U1217 ( .A1(n1173), .A2(n1176), .ZN(n1178) );
  IOA21D1BWP U1218 ( .A1(n1087), .A2(n1040), .B(n1014), .ZN(n1079) );
  OAI222D1BWP U1219 ( .A1(n1116), .A2(n1086), .B1(n1118), .B2(n1078), .C1(n758), .C2(n1013), .ZN(n1087) );
  ND4D1BWP U1220 ( .A1(n1064), .A2(n1038), .A3(n1037), .A4(n1065), .ZN(n1039)
         );
  AOI211XD0BWP U1221 ( .A1(n1071), .A2(n1075), .B(n1072), .C(n1036), .ZN(n1037) );
  OAI21D1BWP U1222 ( .A1(n1055), .A2(n1054), .B(n1068), .ZN(n1036) );
  OAI21D1BWP U1223 ( .A1(n1035), .A2(n1034), .B(n1033), .ZN(n1061) );
  NR2XD0BWP U1224 ( .A1(n1032), .A2(n1116), .ZN(n1035) );
  OAI31D1BWP U1225 ( .A1(n1116), .A2(n1031), .A3(n1030), .B(n1029), .ZN(n1072)
         );
  OAI21D1BWP U1226 ( .A1(n1116), .A2(n1030), .B(n1031), .ZN(n1029) );
  OR2XD1BWP U1227 ( .A1(n1060), .A2(n1026), .Z(n1075) );
  NR2XD0BWP U1228 ( .A1(n1025), .A2(n1024), .ZN(n1071) );
  NR2XD0BWP U1229 ( .A1(n1023), .A2(n1116), .ZN(n1024) );
  XNR2D1BWP U1230 ( .A1(n1060), .A2(n1059), .ZN(n1038) );
  OAI31D1BWP U1231 ( .A1(n1116), .A2(n1022), .A3(n1021), .B(n1020), .ZN(n1026)
         );
  OAI21D1BWP U1232 ( .A1(n1116), .A2(n1021), .B(n1022), .ZN(n1020) );
  IND2D1BWP U1233 ( .A1(n1056), .B1(n1064), .ZN(n1060) );
  INR2D1BWP U1234 ( .A1(n1034), .B1(n1065), .ZN(n1055) );
  AOI21D1BWP U1235 ( .A1(n1019), .A2(n1033), .B(n1018), .ZN(n1054) );
  NR2XD0BWP U1236 ( .A1(n1015), .A2(n1116), .ZN(n1018) );
  OAI222D1BWP U1237 ( .A1(n1118), .A2(n1114), .B1(n1116), .B2(n1117), .C1(
        n1086), .C2(n758), .ZN(n1174) );
  AOI222D1BWP U1238 ( .A1(n1085), .A2(n1084), .B1(n1083), .B2(n1082), .C1(
        n1081), .C2(n759), .ZN(n1117) );
  OAI21D1BWP U1239 ( .A1(n1315), .A2(n1042), .B(n1041), .ZN(n1081) );
  OAI31D1BWP U1240 ( .A1(n1051), .A2(n1000), .A3(n999), .B(n998), .ZN(n1027)
         );
  OAI21D1BWP U1241 ( .A1(n1051), .A2(n999), .B(n1000), .ZN(n998) );
  NR2XD0BWP U1242 ( .A1(n1021), .A2(n1022), .ZN(n1028) );
  NR2XD0BWP U1243 ( .A1(n1016), .A2(n1015), .ZN(n996) );
  IND2D1BWP U1244 ( .A1(n1019), .B1(n1017), .ZN(n1015) );
  NR2XD0BWP U1245 ( .A1(n1032), .A2(n995), .ZN(n1017) );
  XOR2D1BWP U1246 ( .A1(n758), .A2(n994), .Z(n1032) );
  XOR2D1BWP U1247 ( .A1(n993), .A2(n992), .Z(n1016) );
  OAI31D1BWP U1248 ( .A1(n1051), .A2(n991), .A3(n990), .B(n989), .ZN(n997) );
  OAI21D1BWP U1249 ( .A1(n1051), .A2(n990), .B(n991), .ZN(n989) );
  OAI21D1BWP U1250 ( .A1(n988), .A2(n987), .B(n992), .ZN(n1019) );
  AOI21D1BWP U1251 ( .A1(n995), .A2(n985), .B(n987), .ZN(n1034) );
  NR2XD0BWP U1252 ( .A1(n984), .A2(n1051), .ZN(n987) );
  IAO21D1BWP U1253 ( .A1(n1005), .A2(n1078), .B(n1004), .ZN(n1014) );
  OAI222D1BWP U1254 ( .A1(n1118), .A2(n1086), .B1(n1116), .B2(n1114), .C1(
        n1078), .C2(n758), .ZN(n1143) );
  AOI222D1BWP U1255 ( .A1(n1082), .A2(n1012), .B1(n759), .B2(n1077), .C1(n1003), .C2(n1084), .ZN(n1078) );
  AOI222D1BWP U1256 ( .A1(n1077), .A2(n1084), .B1(n1085), .B2(n1082), .C1(
        n1083), .C2(n759), .ZN(n1114) );
  OAI222D1BWP U1257 ( .A1(n1048), .A2(n1047), .B1(n1315), .B2(n1046), .C1(
        n1045), .C2(n766), .ZN(n1083) );
  AOI21D1BWP U1258 ( .A1(n1009), .A2(n1008), .B(n977), .ZN(n1046) );
  AO22D1BWP U1259 ( .A1(n1006), .A2(n1007), .B1(n1314), .B2(n976), .Z(n977) );
  MUX2ND0BWP U1260 ( .I0(n628), .I1(n627), .S(n762), .ZN(n976) );
  AOI222D1BWP U1261 ( .A1(n1012), .A2(n1084), .B1(n1077), .B2(n1082), .C1(
        n1085), .C2(n759), .ZN(n1086) );
  OAI222D1BWP U1262 ( .A1(n1048), .A2(n1045), .B1(n1315), .B2(n1047), .C1(
        n1011), .C2(n766), .ZN(n1085) );
  AOI222D1BWP U1263 ( .A1(n1010), .A2(n1009), .B1(n1008), .B2(n1007), .C1(
        n1006), .C2(n1314), .ZN(n1047) );
  OAI211D1BWP U1264 ( .A1(n626), .A2(n1313), .B(n625), .C(n624), .ZN(n1006) );
  AOI21D1BWP U1265 ( .A1(n684), .A2(N116), .B(n622), .ZN(n625) );
  OAI22D1BWP U1266 ( .A1(n633), .A2(n713), .B1(n709), .B2(n651), .ZN(n622) );
  OAI222D1BWP U1267 ( .A1(n1002), .A2(n766), .B1(n1011), .B2(n1048), .C1(n1045), .C2(n1315), .ZN(n1077) );
  AOI222D1BWP U1268 ( .A1(n1007), .A2(n1010), .B1(n1314), .B2(n1008), .C1(
        n1001), .C2(n1009), .ZN(n1045) );
  OAI21D1BWP U1269 ( .A1(n637), .A2(n691), .B(n636), .ZN(n1008) );
  AOI211XD0BWP U1270 ( .A1(N115), .A2(n761), .B(n635), .C(n634), .ZN(n636) );
  OAI22D1BWP U1271 ( .A1(n633), .A2(n651), .B1(n709), .B2(n657), .ZN(n634) );
  NR2XD0BWP U1272 ( .A1(n713), .A2(n632), .ZN(n635) );
  OAI211D1BWP U1273 ( .A1(n966), .A2(n1025), .B(n1000), .C(n965), .ZN(n967) );
  AOI21D1BWP U1274 ( .A1(n984), .A2(n964), .B(n995), .ZN(n965) );
  OAI21D1BWP U1275 ( .A1(n963), .A2(n962), .B(n961), .ZN(n995) );
  NR2XD0BWP U1276 ( .A1(n960), .A2(n1050), .ZN(n962) );
  OAI31D1BWP U1277 ( .A1(n1050), .A2(n959), .A3(n958), .B(n957), .ZN(n1000) );
  OAI21D1BWP U1278 ( .A1(n1050), .A2(n958), .B(n959), .ZN(n957) );
  NR2XD0BWP U1279 ( .A1(n958), .A2(n953), .ZN(n954) );
  IND2D1BWP U1280 ( .A1(n990), .B1(n991), .ZN(n999) );
  XOR2D1BWP U1281 ( .A1(n990), .A2(n991), .Z(n968) );
  OAI31D1BWP U1282 ( .A1(n1050), .A2(n952), .A3(n951), .B(n950), .ZN(n991) );
  OAI21D1BWP U1283 ( .A1(n1050), .A2(n951), .B(n952), .ZN(n950) );
  NR2XD0BWP U1284 ( .A1(n964), .A2(n984), .ZN(n986) );
  AOI21D1BWP U1285 ( .A1(n948), .A2(n961), .B(n947), .ZN(n988) );
  XOR2D1BWP U1286 ( .A1(n960), .A2(n1050), .Z(n983) );
  XNR2D1BWP U1287 ( .A1(n947), .A2(n945), .ZN(n993) );
  NR2XD0BWP U1288 ( .A1(n944), .A2(n1050), .ZN(n947) );
  OAI21D1BWP U1289 ( .A1(n1013), .A2(n975), .B(n974), .ZN(n1004) );
  AOI222D1BWP U1290 ( .A1(n972), .A2(n1084), .B1(n1003), .B2(n1082), .C1(n1012), .C2(n759), .ZN(n1013) );
  OAI222D1BWP U1291 ( .A1(n1048), .A2(n1002), .B1(n1315), .B2(n1011), .C1(n971), .C2(n766), .ZN(n1012) );
  AOI222D1BWP U1292 ( .A1(n970), .A2(n1009), .B1(n1001), .B2(n1007), .C1(n1010), .C2(n1314), .ZN(n1011) );
  OAI21D1BWP U1293 ( .A1(n713), .A2(n691), .B(n631), .ZN(n1010) );
  AOI211XD0BWP U1294 ( .A1(N116), .A2(n761), .B(n630), .C(n629), .ZN(n631) );
  OAI22D1BWP U1295 ( .A1(n633), .A2(n657), .B1(n709), .B2(n662), .ZN(n629) );
  NR2XD0BWP U1296 ( .A1(n651), .A2(n632), .ZN(n630) );
  NR2XD0BWP U1297 ( .A1(n1084), .A2(n759), .ZN(n1082) );
  OAI22D1BWP U1298 ( .A1(n590), .A2(n589), .B1(n588), .B2(n591), .ZN(N1782) );
  NR2XD0BWP U1299 ( .A1(n1050), .A2(n758), .ZN(n757) );
  AOI21D1BWP U1300 ( .A1(n918), .A2(n1003), .B(n917), .ZN(n974) );
  OAI222D1BWP U1301 ( .A1(n1048), .A2(n971), .B1(n1315), .B2(n1002), .C1(n916), 
        .C2(n766), .ZN(n1003) );
  AOI222D1BWP U1302 ( .A1(n915), .A2(n1009), .B1(n970), .B2(n1007), .C1(n1001), 
        .C2(n1314), .ZN(n1002) );
  OAI21D1BWP U1303 ( .A1(n691), .A2(n651), .B(n621), .ZN(n1001) );
  AOI211XD0BWP U1304 ( .A1(N119), .A2(n684), .B(n620), .C(n619), .ZN(n621) );
  OAI22D1BWP U1305 ( .A1(n633), .A2(n662), .B1(n709), .B2(n667), .ZN(n619) );
  NR2XD0BWP U1306 ( .A1(n713), .A2(n1313), .ZN(n620) );
  NR2XD0BWP U1307 ( .A1(n939), .A2(n938), .ZN(n973) );
  AO211D1BWP U1308 ( .A1(n958), .A2(n956), .B(n953), .C(n935), .Z(n936) );
  IND2D1BWP U1309 ( .A1(n945), .B1(n960), .ZN(n935) );
  OAI31D1BWP U1310 ( .A1(n934), .A2(n933), .A3(n1084), .B(n932), .ZN(n959) );
  OAI21D1BWP U1311 ( .A1(n934), .A2(n1084), .B(n933), .ZN(n932) );
  XNR2D1BWP U1312 ( .A1(n952), .A2(n949), .ZN(n937) );
  NR2XD0BWP U1313 ( .A1(n944), .A2(n945), .ZN(n949) );
  XOR2D1BWP U1314 ( .A1(n930), .A2(n929), .Z(n945) );
  IND2D1BWP U1315 ( .A1(n948), .B1(n946), .ZN(n944) );
  NR2XD0BWP U1316 ( .A1(n960), .A2(n928), .ZN(n946) );
  OAI31D1BWP U1317 ( .A1(n926), .A2(n925), .A3(n1084), .B(n924), .ZN(n952) );
  OAI21D1BWP U1318 ( .A1(n926), .A2(n1084), .B(n925), .ZN(n924) );
  OAI21D1BWP U1319 ( .A1(n923), .A2(n922), .B(n929), .ZN(n948) );
  AOI21D1BWP U1320 ( .A1(n928), .A2(n920), .B(n922), .ZN(n963) );
  INR2D1BWP U1321 ( .A1(n919), .B1(n1084), .ZN(n922) );
  OR2XD1BWP U1322 ( .A1(n927), .A2(n1084), .Z(n920) );
  OAI222D1BWP U1323 ( .A1(n1084), .A2(n1316), .B1(n981), .B2(n943), .C1(n1317), 
        .C2(n980), .ZN(n590) );
  IAO21D1BWP U1324 ( .A1(n1314), .A2(n978), .B(n563), .ZN(n980) );
  AOI222D1BWP U1325 ( .A1(n627), .A2(n914), .B1(n1313), .B2(n626), .C1(n561), 
        .C2(n762), .ZN(n978) );
  AOI21D1BWP U1326 ( .A1(n684), .A2(N115), .B(n560), .ZN(n626) );
  OAI21D1BWP U1327 ( .A1(n913), .A2(n704), .B(n559), .ZN(n560) );
  AOI22D1BWP U1328 ( .A1(n609), .A2(N116), .B1(N127), .B2(N117), .ZN(n559) );
  NR2XD0BWP U1329 ( .A1(n591), .A2(n759), .ZN(n706) );
  IOA21D1BWP U1330 ( .A1(n904), .A2(n903), .B(n902), .ZN(n928) );
  IND2D1BWP U1331 ( .A1(n926), .B1(n925), .ZN(n934) );
  AOI21D1BWP U1332 ( .A1(n896), .A2(n902), .B(n895), .ZN(n923) );
  NR2XD0BWP U1333 ( .A1(n904), .A2(n927), .ZN(n919) );
  OAI31D1BWP U1334 ( .A1(n1315), .A2(n893), .A3(n892), .B(n891), .ZN(n925) );
  OAI21D1BWP U1335 ( .A1(n1315), .A2(n892), .B(n893), .ZN(n891) );
  NR2XD0BWP U1336 ( .A1(n888), .A2(n1315), .ZN(n895) );
  IOA21D1BWP U1337 ( .A1(n972), .A2(n911), .B(n910), .ZN(n917) );
  OAI222D1BWP U1338 ( .A1(n1315), .A2(n971), .B1(n1048), .B2(n916), .C1(n766), 
        .C2(n907), .ZN(n972) );
  AOI222D1BWP U1339 ( .A1(n906), .A2(n1009), .B1(n915), .B2(n1007), .C1(n970), 
        .C2(n1314), .ZN(n971) );
  OAI21D1BWP U1340 ( .A1(n691), .A2(n657), .B(n618), .ZN(n970) );
  AOI211XD0BWP U1341 ( .A1(N120), .A2(n684), .B(n617), .C(n616), .ZN(n618) );
  OAI22D1BWP U1342 ( .A1(n633), .A2(n667), .B1(n709), .B2(n669), .ZN(n616) );
  NR2XD0BWP U1343 ( .A1(n651), .A2(n1313), .ZN(n617) );
  OAI222D1BWP U1344 ( .A1(n1084), .A2(n760), .B1(n1316), .B2(n981), .C1(n943), 
        .C2(n1317), .ZN(n591) );
  AOI21D1BWP U1345 ( .A1(n766), .A2(n570), .B(n558), .ZN(n943) );
  AOI222D1BWP U1346 ( .A1(n627), .A2(n1313), .B1(n557), .B2(n762), .C1(n561), 
        .C2(n914), .ZN(n940) );
  OAI21D1BWP U1347 ( .A1(N114), .A2(n632), .B(n556), .ZN(n627) );
  OA21D1BWP U1348 ( .A1(n941), .A2(n699), .B(n555), .Z(n1316) );
  AOI22D1BWP U1349 ( .A1(n912), .A2(n570), .B1(n698), .B2(n562), .ZN(n555) );
  AO222D1BWP U1350 ( .A1(n554), .A2(n762), .B1(n557), .B2(n914), .C1(n561), 
        .C2(n1313), .Z(n562) );
  OAI222D1BWP U1351 ( .A1(n632), .A2(N113), .B1(n913), .B2(N112), .C1(N114), 
        .C2(n597), .ZN(n561) );
  AOI21D1BWP U1352 ( .A1(n912), .A2(n572), .B(n571), .ZN(n760) );
  AO222D1BWP U1353 ( .A1(n553), .A2(n762), .B1(n554), .B2(n914), .C1(n1313), 
        .C2(n557), .Z(n570) );
  OAI222D1BWP U1354 ( .A1(n632), .A2(N112), .B1(n913), .B2(N111), .C1(N113), 
        .C2(n597), .ZN(n557) );
  AOI211XD0BWP U1355 ( .A1(n914), .A2(n569), .B(n568), .C(n567), .ZN(n697) );
  OAI21D1BWP U1356 ( .A1(N109), .A2(n691), .B(n566), .ZN(n567) );
  NR2XD0BWP U1357 ( .A1(n1009), .A2(n690), .ZN(n568) );
  AOI21D1BWP U1358 ( .A1(n684), .A2(n682), .B(n565), .ZN(n690) );
  OAI22D1BWP U1359 ( .A1(N109), .A2(n597), .B1(N107), .B2(n913), .ZN(n565) );
  AOI222D1BWP U1360 ( .A1(n554), .A2(n1313), .B1(n569), .B2(n762), .C1(n553), 
        .C2(n914), .ZN(n699) );
  NR2XD0BWP U1361 ( .A1(n1313), .A2(n762), .ZN(n914) );
  OAI21D1BWP U1362 ( .A1(N109), .A2(n913), .B(n566), .ZN(n553) );
  AOI22D1BWP U1363 ( .A1(n684), .A2(n688), .B1(n683), .B2(n694), .ZN(n566) );
  OAI21D1BWP U1364 ( .A1(N108), .A2(n913), .B(n689), .ZN(n569) );
  AOI22D1BWP U1365 ( .A1(n684), .A2(n686), .B1(n683), .B2(n688), .ZN(n689) );
  OAI222D1BWP U1366 ( .A1(n632), .A2(N111), .B1(n913), .B2(N110), .C1(N112), 
        .C2(n597), .ZN(n554) );
  IAO21D1BWP U1367 ( .A1(n909), .A2(n916), .B(n908), .ZN(n910) );
  OAI21D1BWP U1368 ( .A1(n907), .A2(n887), .B(n886), .ZN(n908) );
  AOI222D1BWP U1369 ( .A1(n884), .A2(n1009), .B1(n905), .B2(n1007), .C1(n906), 
        .C2(n1314), .ZN(n907) );
  AOI222D1BWP U1370 ( .A1(n1007), .A2(n906), .B1(n1314), .B2(n915), .C1(n905), 
        .C2(n1009), .ZN(n916) );
  OAI21D1BWP U1371 ( .A1(n691), .A2(n662), .B(n615), .ZN(n915) );
  AOI211XD0BWP U1372 ( .A1(N121), .A2(n684), .B(n614), .C(n613), .ZN(n615) );
  OAI22D1BWP U1373 ( .A1(n633), .A2(n669), .B1(n709), .B2(n671), .ZN(n613) );
  NR2XD0BWP U1374 ( .A1(n657), .A2(n1313), .ZN(n614) );
  OAI21D1BWP U1375 ( .A1(n691), .A2(n667), .B(n612), .ZN(n906) );
  AOI211XD0BWP U1376 ( .A1(N122), .A2(n684), .B(n611), .C(n610), .ZN(n612) );
  OAI22D1BWP U1377 ( .A1(n674), .A2(n709), .B1(n633), .B2(n671), .ZN(n610) );
  NR2XD0BWP U1378 ( .A1(n662), .A2(n1313), .ZN(n611) );
  NR2XD0BWP U1379 ( .A1(n1009), .A2(n1314), .ZN(n1007) );
  OAI31D1BWP U1380 ( .A1(n883), .A2(n882), .A3(n941), .B(n881), .ZN(n899) );
  OAI21D1BWP U1381 ( .A1(n883), .A2(n941), .B(n882), .ZN(n881) );
  OAI21D1BWP U1382 ( .A1(n879), .A2(n878), .B(n877), .ZN(n904) );
  NR2XD0BWP U1383 ( .A1(n941), .A2(n876), .ZN(n878) );
  NR2XD0BWP U1384 ( .A1(n888), .A2(n889), .ZN(n890) );
  XOR2D1BWP U1385 ( .A1(n875), .A2(n874), .Z(n889) );
  IND2D1BWP U1386 ( .A1(n896), .B1(n894), .ZN(n888) );
  OAI31D1BWP U1387 ( .A1(n873), .A2(n872), .A3(n941), .B(n871), .ZN(n893) );
  OAI21D1BWP U1388 ( .A1(n873), .A2(n941), .B(n872), .ZN(n871) );
  OAI21D1BWP U1389 ( .A1(n870), .A2(n869), .B(n875), .ZN(n896) );
  AOI21D1BWP U1390 ( .A1(n866), .A2(n905), .B(n865), .ZN(n886) );
  OAI222D1BWP U1391 ( .A1(n667), .A2(n1313), .B1(n752), .B2(n608), .C1(n669), 
        .C2(n691), .ZN(n905) );
  ND4D1BWP U1392 ( .A1(n874), .A2(n862), .A3(n861), .A4(n876), .ZN(n863) );
  AOI211XD0BWP U1393 ( .A1(n860), .A2(n883), .B(n880), .C(n859), .ZN(n861) );
  OAI21D1BWP U1394 ( .A1(n870), .A2(n867), .B(n879), .ZN(n859) );
  OAI31D1BWP U1395 ( .A1(n698), .A2(n855), .A3(n854), .B(n853), .ZN(n880) );
  OAI21D1BWP U1396 ( .A1(n698), .A2(n854), .B(n855), .ZN(n853) );
  IND2D1BWP U1397 ( .A1(n873), .B1(n872), .ZN(n883) );
  XNR2D1BWP U1398 ( .A1(n872), .A2(n873), .ZN(n862) );
  AOI21D1BWP U1399 ( .A1(n852), .A2(n857), .B(n851), .ZN(n870) );
  NR2XD0BWP U1400 ( .A1(n858), .A2(n876), .ZN(n867) );
  OAI31D1BWP U1401 ( .A1(n698), .A2(n849), .A3(n848), .B(n847), .ZN(n872) );
  OAI21D1BWP U1402 ( .A1(n698), .A2(n848), .B(n849), .ZN(n847) );
  XOR2D1BWP U1403 ( .A1(n846), .A2(n851), .Z(n874) );
  IOA21D1BWP U1404 ( .A1(n884), .A2(n844), .B(n763), .ZN(n865) );
  OAI21D1BWP U1405 ( .A1(n608), .A2(n691), .B(n606), .ZN(n884) );
  AOI21D1BWP U1406 ( .A1(n761), .A2(N122), .B(n605), .ZN(n606) );
  OAI21D1BWP U1407 ( .A1(n632), .A2(n674), .B(n604), .ZN(n605) );
  AOI22D1BWP U1408 ( .A1(N125), .A2(n609), .B1(N127), .B2(N126), .ZN(n604) );
  AOI31D1BWP U1409 ( .A1(n843), .A2(n842), .A3(n841), .B(n864), .ZN(n885) );
  ND4D1BWP U1410 ( .A1(n839), .A2(n838), .A3(n837), .A4(n836), .ZN(n840) );
  AOI211XD0BWP U1411 ( .A1(n835), .A2(n607), .B(n833), .C(n834), .ZN(n836) );
  XNR2D1BWP U1412 ( .A1(n830), .A2(n829), .ZN(n838) );
  AOI211XD0BWP U1413 ( .A1(n854), .A2(n607), .B(n828), .C(n855), .ZN(n841) );
  OAI31D1BWP U1414 ( .A1(n835), .A2(n834), .A3(n1009), .B(n827), .ZN(n855) );
  OAI21D1BWP U1415 ( .A1(n835), .A2(n1009), .B(n834), .ZN(n827) );
  IND2D1BWP U1416 ( .A1(n829), .B1(n830), .ZN(n835) );
  IND2D1BWP U1417 ( .A1(n848), .B1(n849), .ZN(n854) );
  XNR2D1BWP U1418 ( .A1(n849), .A2(n848), .ZN(n842) );
  INR2D1BWP U1419 ( .A1(n850), .B1(n852), .ZN(n845) );
  NR2XD0BWP U1420 ( .A1(n856), .A2(n823), .ZN(n850) );
  OAI31D1BWP U1421 ( .A1(n829), .A2(n830), .A3(n1009), .B(n821), .ZN(n849) );
  OAI21D1BWP U1422 ( .A1(n829), .A2(n1009), .B(n830), .ZN(n821) );
  XOR2D1BWP U1423 ( .A1(n818), .A2(n817), .Z(n832) );
  NR2XD0BWP U1424 ( .A1(n858), .A2(n852), .ZN(n843) );
  OAI21D1BWP U1425 ( .A1(n839), .A2(n816), .B(n822), .ZN(n852) );
  NR2XD0BWP U1426 ( .A1(n815), .A2(n814), .ZN(n819) );
  IOA21D1BWP U1427 ( .A1(n813), .A2(n812), .B(n817), .ZN(n814) );
  IND2D1BWP U1428 ( .A1(n811), .B1(n761), .ZN(n817) );
  OAI21D1BWP U1429 ( .A1(n837), .A2(n810), .B(n809), .ZN(n858) );
  NR2XD0BWP U1430 ( .A1(n1009), .A2(n815), .ZN(n816) );
  OR2XD1BWP U1431 ( .A1(n831), .A2(n808), .Z(n815) );
  NR2XD0BWP U1432 ( .A1(n1009), .A2(n831), .ZN(n810) );
  OAI31D1BWP U1433 ( .A1(n804), .A2(n803), .A3(n913), .B(n802), .ZN(n824) );
  OAI21D1BWP U1434 ( .A1(n804), .A2(n913), .B(n803), .ZN(n802) );
  OR2XD1BWP U1435 ( .A1(n801), .A2(n800), .Z(n804) );
  XOR2D1BWP U1436 ( .A1(n826), .A2(n825), .Z(n820) );
  NR2XD0BWP U1437 ( .A1(n818), .A2(n811), .ZN(n825) );
  IND2D1BWP U1438 ( .A1(n813), .B1(n799), .ZN(n811) );
  OAI21D1BWP U1439 ( .A1(n798), .A2(n797), .B(n796), .ZN(n813) );
  XOR2D1BWP U1440 ( .A1(n796), .A2(n795), .Z(n818) );
  OAI31D1BWP U1441 ( .A1(n801), .A2(n793), .A3(n913), .B(n792), .ZN(n826) );
  OAI21D1BWP U1442 ( .A1(n801), .A2(n913), .B(n793), .ZN(n792) );
  OA21D1BWP U1443 ( .A1(n608), .A2(n806), .B(n552), .Z(n763) );
  AOI222D1BWP U1444 ( .A1(N125), .A2(N127), .B1(n597), .B2(N123), .C1(N124), 
        .C2(n609), .ZN(n608) );
  NR2XD0BWP U1445 ( .A1(N127), .A2(n597), .ZN(n609) );
  IOA21D1BWP U1446 ( .A1(n808), .A2(n791), .B(n812), .ZN(n823) );
  INR2D1BWP U1447 ( .A1(n807), .B1(n790), .ZN(n799) );
  AOI21D1BWP U1448 ( .A1(n551), .A2(N124), .B(n550), .ZN(n552) );
  AO21D1BWP U1449 ( .A1(n603), .A2(n602), .B(n601), .Z(n800) );
  NR2XD0BWP U1450 ( .A1(n788), .A2(n787), .ZN(n794) );
  OR2XD1BWP U1451 ( .A1(n600), .A2(n601), .Z(n803) );
  NR2XD0BWP U1452 ( .A1(n602), .A2(n603), .ZN(n601) );
  OAI21D1BWP U1453 ( .A1(n753), .A2(n785), .B(n786), .ZN(n788) );
  ND4D1BWP U1454 ( .A1(n753), .A2(n597), .A3(n596), .A4(n595), .ZN(n786) );
  AO21D1BWP U1455 ( .A1(n790), .A2(n784), .B(n797), .Z(n808) );
  NR2XD0BWP U1456 ( .A1(n913), .A2(n787), .ZN(n797) );
  XNR2D1BWP U1457 ( .A1(n592), .A2(n597), .ZN(n789) );
  MUX2ND0BWP U1458 ( .I0(n779), .I1(n1344), .S(N127), .ZN(n599) );
  MUX2ND0BWP U1459 ( .I0(n781), .I1(n642), .S(N127), .ZN(n600) );
  OAI22D1BWP U1460 ( .A1(N127), .A2(n777), .B1(n776), .B2(B[14]), .ZN(n607) );
  NR2XD0BWP U1461 ( .A1(n775), .A2(n1343), .ZN(n780) );
  MUX2ND0BWP U1462 ( .I0(n1334), .I1(n1333), .S(n548), .ZN(n753) );
  MUX2ND0BWP U1463 ( .I0(n1308), .I1(n1343), .S(n547), .ZN(n603) );
  NR2XD0BWP U1464 ( .A1(N127), .A2(n775), .ZN(n547) );
  IND2D1BWP U1465 ( .A1(n778), .B1(n1341), .ZN(n775) );
  NR2XD0BWP U1466 ( .A1(n594), .A2(n593), .ZN(n785) );
  MUX2ND0BWP U1467 ( .I0(n1326), .I1(n1337), .S(N127), .ZN(n592) );
  AOI21D1BWP U1468 ( .A1(n1344), .A2(n778), .B(n773), .ZN(n782) );
  OAI211D1BWP U1469 ( .A1(n1344), .A2(n778), .B(n1238), .C(n772), .ZN(n773) );
  MUX2D1BWP U1470 ( .I0(n1329), .I1(n1328), .S(N127), .Z(n596) );
  NR2XD0BWP U1471 ( .A1(n1326), .A2(n1335), .ZN(n774) );
  ND4D1BWP U1472 ( .A1(B[11]), .A2(B[13]), .A3(B[12]), .A4(n1321), .ZN(n1346)
         );
  NR2XD0BWP U1473 ( .A1(n764), .A2(n765), .ZN(n1321) );
  OAI21D1BWP U1474 ( .A1(n1338), .A2(n1239), .B(n1238), .ZN(n1323) );
  INVD1BWP U1475 ( .I(B[9]), .ZN(n534) );
  NR2XD0BWP U1476 ( .A1(B[14]), .A2(n776), .ZN(n1310) );
  TIELBWP U1477 ( .ZN(operprod[22]) );
  FA1D0BWP U1478 ( .A(A[11]), .B(B[11]), .CI(n768), .CO(n769), .S(n1335) );
  FA1D0BWP U1479 ( .A(A[12]), .B(B[12]), .CI(n769), .CO(n770), .S(n1333) );
  FA1D0BWP U1480 ( .A(n764), .B(A[14]), .CI(n771), .CO(n776), .S(n1343) );
  NR4D0BWP U1481 ( .A1(n1337), .A2(n1333), .A3(n1335), .A4(n1343), .ZN(n772)
         );
  MUX2ND0BWP U1482 ( .I0(n1344), .I1(n1341), .S(n778), .ZN(n779) );
  MUX2ND0BWP U1483 ( .I0(n1238), .I1(n642), .S(n780), .ZN(n781) );
  MUX2ND0BWP U1484 ( .I0(n913), .I1(n752), .S(n789), .ZN(n807) );
  NR4D0BWP U1485 ( .A1(n807), .A2(n813), .A3(n818), .A4(n808), .ZN(n805) );
  MUX2ND0BWP U1486 ( .I0(n761), .I1(n1313), .S(n807), .ZN(n831) );
  INR4D0BWP U1487 ( .A1(n963), .B1(n948), .B2(n937), .B3(n936), .ZN(n938) );
  MUX2ND0BWP U1488 ( .I0(n979), .I1(n978), .S(n766), .ZN(n1042) );
  OA22D1BWP U1489 ( .A1(n1048), .A2(n1046), .B1(n766), .B2(n1047), .Z(n1041)
         );
  MUX2ND0BWP U1490 ( .I0(n1081), .I1(n1043), .S(n1319), .ZN(n1049) );
  MUX2ND0BWP U1491 ( .I0(n1113), .I1(n1175), .S(n1173), .ZN(n1120) );
  INR4D0BWP U1492 ( .A1(n1167), .B1(n1151), .B2(n1140), .B3(n1139), .ZN(n1142)
         );
  MUX2ND0BWP U1493 ( .I0(n1144), .I1(n1179), .S(n1181), .ZN(n1180) );
  NR4D0BWP U1494 ( .A1(n1201), .A2(n1206), .A3(n1172), .A4(n1171), .ZN(n1209)
         );
  MUX2ND0BWP U1495 ( .I0(n1179), .I1(n1183), .S(n1181), .ZN(n1186) );
  MUX2ND0BWP U1496 ( .I0(n1183), .I1(n1182), .S(n1181), .ZN(n1185) );
  MUX2ND0BWP U1497 ( .I0(n1186), .I1(n1185), .S(n1184), .ZN(n1187) );
  MUX2ND0BWP U1498 ( .I0(n754), .I1(n1187), .S(n755), .ZN(n1210) );
  NR3D0BWP U1499 ( .A1(n1337), .A2(n1334), .A3(n1239), .ZN(n1237) );
  INR3D0BWP U1500 ( .A1(n1306), .B1(n1280), .B2(n1284), .ZN(n1277) );
  INR4D0BWP U1501 ( .A1(n1330), .B1(n1307), .B2(n1309), .B3(n1302), .ZN(n1304)
         );
endmodule



    