module DRAM(output [15:0] DataOut, input [15:0] Addr, input Clk1, input Clk2,
    input [15:0] DataIn, input RD, input WR);
    
endmodule
