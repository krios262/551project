module VADD16(output [255:0] SumV,output Overflw,input [255:0] Inval1,input [255:0] Inval2,input start,output done);

  wire [15:0] Ov;

  assign Overflw = Ov[0] |Ov[1] | Ov[2] | Ov[3] | Ov[4] | Ov[5] | Ov[6] | Ov[7] | Ov[8] | Ov[9] | Ov[10] | Ov[11] | Ov[12] | Ov[13] | Ov[14] | Ov[15] ; 
  assign done = start;

  VADD adder[15:0](SumV,Ov,Inval1,Inval2);
  /*
  VADD add1(SumV[15:0],Ov[0],Inval1[15:0],Inval2[15:0]);
  VADD add2(SumV[31:16],Ov[1],Inval1[31:16],Inval2[31:16]);
  VADD add3(SumV[47:32],Ov[2],Inval1[47:32],Inval2[47:32]);
  VADD add4(SumV[63:48],Ov[3],Inval1[63:48],Inval2[63:48]);
  VADD add5(SumV[79:64],Ov[4],Inval1[79:64],Inval2[79:64]);
  VADD add6(SumV[95:80],Ov[5],Inval1[95:80],Inval2[95:80]);
  VADD add7(SumV[111:96],Ov[6],Inval1[111:96],Inval2[111:96]);
  VADD add8(SumV[127:112],Ov[7],Inval1[127:112],Inval2[127:112]);
  VADD add9(SumV[143:128],Ov[8],Inval1[143:128],Inval2[143:128]);
  VADD add10(SumV[159:144],Ov[9],Inval1[159:144],Inval2[159:144]);
  VADD add11(SumV[175:160],Ov[10],Inval1[175:160],Inval2[175:160]);
  VADD add12(SumV[191:176],Ov[11],Inval1[191:176],Inval2[191:176]);
  VADD add13(SumV[207:192],Ov[12],Inval1[207:192],Inval2[207:192]);
  VADD add14(SumV[223:208],Ov[13],Inval1[223:208],Inval2[223:208]);
  VADD add15(SumV[239:224],Ov[14],Inval1[239:224],Inval2[239:224]);
  VADD add16(SumV[255:240],Ov[15],Inval1[255:240],Inval2[255:240]);
  */

endmodule
